LIBRARY ieee;
USE ieee.std_logic_textio.ALL;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY effMastrovito IS
	PORT (
		clk : IN STD_LOGIC;
		in_val : IN STD_LOGIC;
		X : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		Y : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		out_val : OUT STD_LOGIC;
		out_product : OUT STD_LOGIC_VECTOR(127 DOWNTO 0));
END ENTITY;

ARCHITECTURE effMastrovito_arc OF effMastrovito IS

	SIGNAL A,B,C : STD_LOGIC_VECTOR(127 DOWNTO 0);
	
BEGIN    

		PROCESS (clk)
		BEGIN
			IF (RISING_EDGE(clk)) THEN
				A <= X;
				B <= Y;
			END IF;
		END PROCESS;
	
    C(0)   <= (A(0) and B(0)) xor (A(0) and B(127)) xor (A(1) and B(126)) xor (A(2) and B(125)) xor (A(3) and B(124)) xor (A(4) and B(123)) xor (A(5) and B(122)) xor (A(6) and B(121)) xor (A(7) and B(120)) xor (A(8) and B(119)) xor (A(9) and B(118)) xor (A(10) and B(117)) xor (A(11) and B(116)) xor (A(12) and B(115)) xor (A(13) and B(114)) xor (A(14) and B(113)) xor (A(15) and B(112)) xor (A(16) and B(111)) xor (A(17) and B(110)) xor (A(18) and B(109)) xor (A(19) and B(108)) xor (A(20) and B(107)) xor (A(21) and B(106)) xor (A(23) and B(105)) xor (A(23) and B(104)) xor (A(24) and B(103)) xor (A(25) and B(102)) xor (A(26) and B(101)) xor (A(27) and B(100)) xor (A(28) and B(99)) xor (A(29) and B(98)) xor (A(30) and B(97)) xor (A(31) and B(96)) xor (A(32) and B(95)) xor (A(33) and B(94)) xor (A(34) and B(93)) xor (A(35) and B(92)) xor (A(36) and B(91)) xor (A(37) and B(90)) xor (A(38) and B(89)) xor (A(39) and B(88)) xor (A(40) and B(87)) xor (A(41) and B(86)) xor (A(42) and B(85)) xor (A(43) and B(84)) xor (A(44) and B(83)) xor (A(45) and B(82)) xor (A(46) and B(81)) xor (A(47) and B(80)) xor (A(48) and B(79)) xor (A(49) and B(78)) xor (A(50) and B(77)) xor (A(51) and B(76)) xor (A(52) and B(75)) xor (A(53) and B(74)) xor (A(54) and B(73)) xor (A(55) and B(72)) xor (A(56) and B(71)) xor (A(57) and B(70)) xor (A(58) and B(69)) xor (A(59) and B(68)) xor (A(60) and B(67)) xor (A(61) and B(66)) xor (A(62) and B(65)) xor (A(63) and B(64)) xor (A(64) and B(63)) xor (A(65) and B(62)) xor (A(66) and B(61)) xor (A(67) and B(60)) xor (A(68) and B(59)) xor (A(69) and B(58)) xor (A(70) and B(57)) xor (A(71) and B(56)) xor (A(72) and B(55)) xor (A(73) and B(54)) xor (A(74) and B(53)) xor (A(75) and B(52)) xor (A(76) and B(51)) xor (A(77) and B(50)) xor (A(78) and B(49)) xor (A(79) and B(48)) xor (A(80) and B(47)) xor (A(81) and B(46)) xor (A(82) and B(45)) xor (A(83) and B(44)) xor (A(84) and B(43)) xor (A(85) and B(42)) xor (A(86) and B(41)) xor (A(87) and B(40)) xor (A(88) and B(39)) xor (A(89) and B(38)) xor (A(90) and B(37)) xor (A(91) and B(36)) xor (A(92) and B(35)) xor (A(93) and B(34)) xor (A(94) and B(33)) xor (A(95) and B(32)) xor (A(96) and B(31)) xor (A(97) and B(30)) xor (A(98) and B(29)) xor (A(99) and B(28)) xor (A(100) and B(27)) xor (A(101) and B(26)) xor (A(102) and B(25)) xor (A(103) and B(24)) xor (A(104) and B(23)) xor (A(105) and B(23)) xor (A(106) and B(21)) xor (A(107) and B(20)) xor (A(108) and B(19)) xor (A(109) and B(18)) xor (A(110) and B(17)) xor (A(111) and B(16)) xor (A(112) and B(15)) xor (A(113) and B(14)) xor (A(114) and B(13)) xor (A(115) and B(12)) xor (A(116) and B(11)) xor (A(117) and B(10)) xor (A(118) and B(9)) xor (A(119) and B(8)) xor (A(120) and B(7)) xor (A(121) and B(6)) xor (A(122) and B(5)) xor (A(123) and B(4)) xor (A(124) and B(3)) xor (A(125) and B(2)) xor (A(126) and B(1)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(122)) xor (A(126) and B(127));
    C(1)   <= (A(0) and B(1)) xor (A(1) and B(0)) xor (A(0) and B(127)) xor (A(1) and B(126)) xor (A(2) and B(125)) xor (A(3) and B(124)) xor (A(4) and B(123)) xor (A(5) and B(122)) xor (A(6) and B(121)) xor (A(7) and B(120)) xor (A(8) and B(119)) xor (A(9) and B(118)) xor (A(10) and B(117)) xor (A(11) and B(116)) xor (A(12) and B(115)) xor (A(13) and B(114)) xor (A(14) and B(113)) xor (A(15) and B(112)) xor (A(16) and B(111)) xor (A(17) and B(110)) xor (A(18) and B(109)) xor (A(19) and B(108)) xor (A(20) and B(107)) xor (A(21) and B(106)) xor (A(23) and B(105)) xor (A(23) and B(104)) xor (A(24) and B(103)) xor (A(25) and B(102)) xor (A(26) and B(101)) xor (A(27) and B(100)) xor (A(28) and B(99)) xor (A(29) and B(98)) xor (A(30) and B(97)) xor (A(31) and B(96)) xor (A(32) and B(95)) xor (A(33) and B(94)) xor (A(34) and B(93)) xor (A(35) and B(92)) xor (A(36) and B(91)) xor (A(37) and B(90)) xor (A(38) and B(89)) xor (A(39) and B(88)) xor (A(40) and B(87)) xor (A(41) and B(86)) xor (A(42) and B(85)) xor (A(43) and B(84)) xor (A(44) and B(83)) xor (A(45) and B(82)) xor (A(46) and B(81)) xor (A(47) and B(80)) xor (A(48) and B(79)) xor (A(49) and B(78)) xor (A(50) and B(77)) xor (A(51) and B(76)) xor (A(52) and B(75)) xor (A(53) and B(74)) xor (A(54) and B(73)) xor (A(55) and B(72)) xor (A(56) and B(71)) xor (A(57) and B(70)) xor (A(58) and B(69)) xor (A(59) and B(68)) xor (A(60) and B(67)) xor (A(61) and B(66)) xor (A(62) and B(65)) xor (A(63) and B(64)) xor (A(64) and B(63)) xor (A(65) and B(62)) xor (A(66) and B(61)) xor (A(67) and B(60)) xor (A(68) and B(59)) xor (A(69) and B(58)) xor (A(70) and B(57)) xor (A(71) and B(56)) xor (A(72) and B(55)) xor (A(73) and B(54)) xor (A(74) and B(53)) xor (A(75) and B(52)) xor (A(76) and B(51)) xor (A(77) and B(50)) xor (A(78) and B(49)) xor (A(79) and B(48)) xor (A(80) and B(47)) xor (A(81) and B(46)) xor (A(82) and B(45)) xor (A(83) and B(44)) xor (A(84) and B(43)) xor (A(85) and B(42)) xor (A(86) and B(41)) xor (A(87) and B(40)) xor (A(88) and B(39)) xor (A(89) and B(38)) xor (A(90) and B(37)) xor (A(91) and B(36)) xor (A(92) and B(35)) xor (A(93) and B(34)) xor (A(94) and B(33)) xor (A(95) and B(32)) xor (A(96) and B(31)) xor (A(97) and B(30)) xor (A(98) and B(29)) xor (A(99) and B(28)) xor (A(100) and B(27)) xor (A(101) and B(26)) xor (A(102) and B(25)) xor (A(103) and B(24)) xor (A(104) and B(23)) xor (A(105) and B(23)) xor (A(106) and B(21)) xor (A(107) and B(20)) xor (A(108) and B(19)) xor (A(109) and B(18)) xor (A(110) and B(17)) xor (A(111) and B(16)) xor (A(112) and B(15)) xor (A(113) and B(14)) xor (A(114) and B(13)) xor (A(115) and B(12)) xor (A(116) and B(11)) xor (A(117) and B(10)) xor (A(118) and B(9)) xor (A(119) and B(8)) xor (A(120) and B(7)) xor (A(121) and B(6)) xor (A(122) and B(5)) xor (A(123) and B(4)) xor (A(124) and B(3)) xor (A(125) and B(2)) xor (A(126) and B(1)) xor (A(1) and B(127)) xor (A(2) and B(126)) xor (A(3) and B(125)) xor (A(4) and B(124)) xor (A(5) and B(123)) xor (A(6) and B(122)) xor (A(7) and B(121)) xor (A(8) and B(120)) xor (A(9) and B(119)) xor (A(10) and B(118)) xor (A(11) and B(117)) xor (A(12) and B(116)) xor (A(13) and B(115)) xor (A(14) and B(114)) xor (A(15) and B(113)) xor (A(16) and B(112)) xor (A(17) and B(111)) xor (A(18) and B(110)) xor (A(19) and B(109)) xor (A(20) and B(108)) xor (A(21) and B(107)) xor (A(23) and B(106)) xor (A(23) and B(105)) xor (A(24) and B(104)) xor (A(25) and B(103)) xor (A(26) and B(102)) xor (A(27) and B(101)) xor (A(28) and B(100)) xor (A(29) and B(99)) xor (A(30) and B(98)) xor (A(31) and B(97)) xor (A(32) and B(96)) xor (A(33) and B(95)) xor (A(34) and B(94)) xor (A(35) and B(93)) xor (A(36) and B(92)) xor (A(37) and B(91)) xor (A(38) and B(90)) xor (A(39) and B(89)) xor (A(40) and B(88)) xor (A(41) and B(87)) xor (A(42) and B(86)) xor (A(43) and B(85)) xor (A(44) and B(84)) xor (A(45) and B(83)) xor (A(46) and B(82)) xor (A(47) and B(81)) xor (A(48) and B(80)) xor (A(49) and B(79)) xor (A(50) and B(78)) xor (A(51) and B(77)) xor (A(52) and B(76)) xor (A(53) and B(75)) xor (A(54) and B(74)) xor (A(55) and B(73)) xor (A(56) and B(72)) xor (A(57) and B(71)) xor (A(58) and B(70)) xor (A(59) and B(69)) xor (A(60) and B(68)) xor (A(61) and B(67)) xor (A(62) and B(66)) xor (A(63) and B(65)) xor (A(64) and B(64)) xor (A(65) and B(63)) xor (A(66) and B(62)) xor (A(67) and B(61)) xor (A(68) and B(60)) xor (A(69) and B(59)) xor (A(70) and B(58)) xor (A(71) and B(57)) xor (A(72) and B(56)) xor (A(73) and B(55)) xor (A(74) and B(54)) xor (A(75) and B(53)) xor (A(76) and B(52)) xor (A(77) and B(51)) xor (A(78) and B(50)) xor (A(79) and B(49)) xor (A(80) and B(48)) xor (A(81) and B(47)) xor (A(82) and B(46)) xor (A(83) and B(45)) xor (A(84) and B(44)) xor (A(85) and B(43)) xor (A(86) and B(42)) xor (A(87) and B(41)) xor (A(88) and B(40)) xor (A(89) and B(39)) xor (A(90) and B(38)) xor (A(91) and B(37)) xor (A(92) and B(36)) xor (A(93) and B(35)) xor (A(94) and B(34)) xor (A(95) and B(33)) xor (A(96) and B(32)) xor (A(97) and B(31)) xor (A(98) and B(30)) xor (A(99) and B(29)) xor (A(100) and B(28)) xor (A(101) and B(27)) xor (A(102) and B(26)) xor (A(103) and B(25)) xor (A(104) and B(24)) xor (A(105) and B(23)) xor (A(106) and B(23)) xor (A(107) and B(21)) xor (A(108) and B(20)) xor (A(109) and B(19)) xor (A(110) and B(18)) xor (A(111) and B(17)) xor (A(112) and B(16)) xor (A(113) and B(15)) xor (A(114) and B(14)) xor (A(115) and B(13)) xor (A(116) and B(12)) xor (A(117) and B(11)) xor (A(118) and B(10)) xor (A(119) and B(9)) xor (A(120) and B(8)) xor (A(121) and B(7)) xor (A(122) and B(6)) xor (A(123) and B(5)) xor (A(124) and B(4)) xor (A(125) and B(3)) xor (A(126) and B(2)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(122)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(123)) xor (A(126) and B(127));
    C(2)   <= (A(0) and B(2)) xor (A(1) and B(1)) xor (A(2) and B(0)) xor (A(0) and B(127)) xor (A(1) and B(126)) xor (A(2) and B(125)) xor (A(3) and B(124)) xor (A(4) and B(123)) xor (A(5) and B(122)) xor (A(6) and B(121)) xor (A(7) and B(120)) xor (A(8) and B(119)) xor (A(9) and B(118)) xor (A(10) and B(117)) xor (A(11) and B(116)) xor (A(12) and B(115)) xor (A(13) and B(114)) xor (A(14) and B(113)) xor (A(15) and B(112)) xor (A(16) and B(111)) xor (A(17) and B(110)) xor (A(18) and B(109)) xor (A(19) and B(108)) xor (A(20) and B(107)) xor (A(21) and B(106)) xor (A(23) and B(105)) xor (A(23) and B(104)) xor (A(24) and B(103)) xor (A(25) and B(102)) xor (A(26) and B(101)) xor (A(27) and B(100)) xor (A(28) and B(99)) xor (A(29) and B(98)) xor (A(30) and B(97)) xor (A(31) and B(96)) xor (A(32) and B(95)) xor (A(33) and B(94)) xor (A(34) and B(93)) xor (A(35) and B(92)) xor (A(36) and B(91)) xor (A(37) and B(90)) xor (A(38) and B(89)) xor (A(39) and B(88)) xor (A(40) and B(87)) xor (A(41) and B(86)) xor (A(42) and B(85)) xor (A(43) and B(84)) xor (A(44) and B(83)) xor (A(45) and B(82)) xor (A(46) and B(81)) xor (A(47) and B(80)) xor (A(48) and B(79)) xor (A(49) and B(78)) xor (A(50) and B(77)) xor (A(51) and B(76)) xor (A(52) and B(75)) xor (A(53) and B(74)) xor (A(54) and B(73)) xor (A(55) and B(72)) xor (A(56) and B(71)) xor (A(57) and B(70)) xor (A(58) and B(69)) xor (A(59) and B(68)) xor (A(60) and B(67)) xor (A(61) and B(66)) xor (A(62) and B(65)) xor (A(63) and B(64)) xor (A(64) and B(63)) xor (A(65) and B(62)) xor (A(66) and B(61)) xor (A(67) and B(60)) xor (A(68) and B(59)) xor (A(69) and B(58)) xor (A(70) and B(57)) xor (A(71) and B(56)) xor (A(72) and B(55)) xor (A(73) and B(54)) xor (A(74) and B(53)) xor (A(75) and B(52)) xor (A(76) and B(51)) xor (A(77) and B(50)) xor (A(78) and B(49)) xor (A(79) and B(48)) xor (A(80) and B(47)) xor (A(81) and B(46)) xor (A(82) and B(45)) xor (A(83) and B(44)) xor (A(84) and B(43)) xor (A(85) and B(42)) xor (A(86) and B(41)) xor (A(87) and B(40)) xor (A(88) and B(39)) xor (A(89) and B(38)) xor (A(90) and B(37)) xor (A(91) and B(36)) xor (A(92) and B(35)) xor (A(93) and B(34)) xor (A(94) and B(33)) xor (A(95) and B(32)) xor (A(96) and B(31)) xor (A(97) and B(30)) xor (A(98) and B(29)) xor (A(99) and B(28)) xor (A(100) and B(27)) xor (A(101) and B(26)) xor (A(102) and B(25)) xor (A(103) and B(24)) xor (A(104) and B(23)) xor (A(105) and B(23)) xor (A(106) and B(21)) xor (A(107) and B(20)) xor (A(108) and B(19)) xor (A(109) and B(18)) xor (A(110) and B(17)) xor (A(111) and B(16)) xor (A(112) and B(15)) xor (A(113) and B(14)) xor (A(114) and B(13)) xor (A(115) and B(12)) xor (A(116) and B(11)) xor (A(117) and B(10)) xor (A(118) and B(9)) xor (A(119) and B(8)) xor (A(120) and B(7)) xor (A(121) and B(6)) xor (A(122) and B(5)) xor (A(123) and B(4)) xor (A(124) and B(3)) xor (A(125) and B(2)) xor (A(126) and B(1)) xor (A(1) and B(127)) xor (A(2) and B(126)) xor (A(3) and B(125)) xor (A(4) and B(124)) xor (A(5) and B(123)) xor (A(6) and B(122)) xor (A(7) and B(121)) xor (A(8) and B(120)) xor (A(9) and B(119)) xor (A(10) and B(118)) xor (A(11) and B(117)) xor (A(12) and B(116)) xor (A(13) and B(115)) xor (A(14) and B(114)) xor (A(15) and B(113)) xor (A(16) and B(112)) xor (A(17) and B(111)) xor (A(18) and B(110)) xor (A(19) and B(109)) xor (A(20) and B(108)) xor (A(21) and B(107)) xor (A(23) and B(106)) xor (A(23) and B(105)) xor (A(24) and B(104)) xor (A(25) and B(103)) xor (A(26) and B(102)) xor (A(27) and B(101)) xor (A(28) and B(100)) xor (A(29) and B(99)) xor (A(30) and B(98)) xor (A(31) and B(97)) xor (A(32) and B(96)) xor (A(33) and B(95)) xor (A(34) and B(94)) xor (A(35) and B(93)) xor (A(36) and B(92)) xor (A(37) and B(91)) xor (A(38) and B(90)) xor (A(39) and B(89)) xor (A(40) and B(88)) xor (A(41) and B(87)) xor (A(42) and B(86)) xor (A(43) and B(85)) xor (A(44) and B(84)) xor (A(45) and B(83)) xor (A(46) and B(82)) xor (A(47) and B(81)) xor (A(48) and B(80)) xor (A(49) and B(79)) xor (A(50) and B(78)) xor (A(51) and B(77)) xor (A(52) and B(76)) xor (A(53) and B(75)) xor (A(54) and B(74)) xor (A(55) and B(73)) xor (A(56) and B(72)) xor (A(57) and B(71)) xor (A(58) and B(70)) xor (A(59) and B(69)) xor (A(60) and B(68)) xor (A(61) and B(67)) xor (A(62) and B(66)) xor (A(63) and B(65)) xor (A(64) and B(64)) xor (A(65) and B(63)) xor (A(66) and B(62)) xor (A(67) and B(61)) xor (A(68) and B(60)) xor (A(69) and B(59)) xor (A(70) and B(58)) xor (A(71) and B(57)) xor (A(72) and B(56)) xor (A(73) and B(55)) xor (A(74) and B(54)) xor (A(75) and B(53)) xor (A(76) and B(52)) xor (A(77) and B(51)) xor (A(78) and B(50)) xor (A(79) and B(49)) xor (A(80) and B(48)) xor (A(81) and B(47)) xor (A(82) and B(46)) xor (A(83) and B(45)) xor (A(84) and B(44)) xor (A(85) and B(43)) xor (A(86) and B(42)) xor (A(87) and B(41)) xor (A(88) and B(40)) xor (A(89) and B(39)) xor (A(90) and B(38)) xor (A(91) and B(37)) xor (A(92) and B(36)) xor (A(93) and B(35)) xor (A(94) and B(34)) xor (A(95) and B(33)) xor (A(96) and B(32)) xor (A(97) and B(31)) xor (A(98) and B(30)) xor (A(99) and B(29)) xor (A(100) and B(28)) xor (A(101) and B(27)) xor (A(102) and B(26)) xor (A(103) and B(25)) xor (A(104) and B(24)) xor (A(105) and B(23)) xor (A(106) and B(23)) xor (A(107) and B(21)) xor (A(108) and B(20)) xor (A(109) and B(19)) xor (A(110) and B(18)) xor (A(111) and B(17)) xor (A(112) and B(16)) xor (A(113) and B(15)) xor (A(114) and B(14)) xor (A(115) and B(13)) xor (A(116) and B(12)) xor (A(117) and B(11)) xor (A(118) and B(10)) xor (A(119) and B(9)) xor (A(120) and B(8)) xor (A(121) and B(7)) xor (A(122) and B(6)) xor (A(123) and B(5)) xor (A(124) and B(4)) xor (A(125) and B(3)) xor (A(126) and B(2)) xor (A(2) and B(127)) xor (A(3) and B(126)) xor (A(4) and B(125)) xor (A(5) and B(124)) xor (A(6) and B(123)) xor (A(7) and B(122)) xor (A(8) and B(121)) xor (A(9) and B(120)) xor (A(10) and B(119)) xor (A(11) and B(118)) xor (A(12) and B(117)) xor (A(13) and B(116)) xor (A(14) and B(115)) xor (A(15) and B(114)) xor (A(16) and B(113)) xor (A(17) and B(112)) xor (A(18) and B(111)) xor (A(19) and B(110)) xor (A(20) and B(109)) xor (A(21) and B(108)) xor (A(23) and B(107)) xor (A(23) and B(106)) xor (A(24) and B(105)) xor (A(25) and B(104)) xor (A(26) and B(103)) xor (A(27) and B(102)) xor (A(28) and B(101)) xor (A(29) and B(100)) xor (A(30) and B(99)) xor (A(31) and B(98)) xor (A(32) and B(97)) xor (A(33) and B(96)) xor (A(34) and B(95)) xor (A(35) and B(94)) xor (A(36) and B(93)) xor (A(37) and B(92)) xor (A(38) and B(91)) xor (A(39) and B(90)) xor (A(40) and B(89)) xor (A(41) and B(88)) xor (A(42) and B(87)) xor (A(43) and B(86)) xor (A(44) and B(85)) xor (A(45) and B(84)) xor (A(46) and B(83)) xor (A(47) and B(82)) xor (A(48) and B(81)) xor (A(49) and B(80)) xor (A(50) and B(79)) xor (A(51) and B(78)) xor (A(52) and B(77)) xor (A(53) and B(76)) xor (A(54) and B(75)) xor (A(55) and B(74)) xor (A(56) and B(73)) xor (A(57) and B(72)) xor (A(58) and B(71)) xor (A(59) and B(70)) xor (A(60) and B(69)) xor (A(61) and B(68)) xor (A(62) and B(67)) xor (A(63) and B(66)) xor (A(64) and B(65)) xor (A(65) and B(64)) xor (A(66) and B(63)) xor (A(67) and B(62)) xor (A(68) and B(61)) xor (A(69) and B(60)) xor (A(70) and B(59)) xor (A(71) and B(58)) xor (A(72) and B(57)) xor (A(73) and B(56)) xor (A(74) and B(55)) xor (A(75) and B(54)) xor (A(76) and B(53)) xor (A(77) and B(52)) xor (A(78) and B(51)) xor (A(79) and B(50)) xor (A(80) and B(49)) xor (A(81) and B(48)) xor (A(82) and B(47)) xor (A(83) and B(46)) xor (A(84) and B(45)) xor (A(85) and B(44)) xor (A(86) and B(43)) xor (A(87) and B(42)) xor (A(88) and B(41)) xor (A(89) and B(40)) xor (A(90) and B(39)) xor (A(91) and B(38)) xor (A(92) and B(37)) xor (A(93) and B(36)) xor (A(94) and B(35)) xor (A(95) and B(34)) xor (A(96) and B(33)) xor (A(97) and B(32)) xor (A(98) and B(31)) xor (A(99) and B(30)) xor (A(100) and B(29)) xor (A(101) and B(28)) xor (A(102) and B(27)) xor (A(103) and B(26)) xor (A(104) and B(25)) xor (A(105) and B(24)) xor (A(106) and B(23)) xor (A(107) and B(23)) xor (A(108) and B(21)) xor (A(109) and B(20)) xor (A(110) and B(19)) xor (A(111) and B(18)) xor (A(112) and B(17)) xor (A(113) and B(16)) xor (A(114) and B(15)) xor (A(115) and B(14)) xor (A(116) and B(13)) xor (A(117) and B(12)) xor (A(118) and B(11)) xor (A(119) and B(10)) xor (A(120) and B(9)) xor (A(121) and B(8)) xor (A(122) and B(7)) xor (A(123) and B(6)) xor (A(124) and B(5)) xor (A(125) and B(4)) xor (A(126) and B(3)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(122)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(123)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(124)) xor (A(126) and B(127));
    C(3)   <= (A(0) and B(3)) xor (A(1) and B(2)) xor (A(2) and B(1)) xor (A(3) and B(0)) xor (A(1) and B(127)) xor (A(2) and B(126)) xor (A(3) and B(125)) xor (A(4) and B(124)) xor (A(5) and B(123)) xor (A(6) and B(122)) xor (A(7) and B(121)) xor (A(8) and B(120)) xor (A(9) and B(119)) xor (A(10) and B(118)) xor (A(11) and B(117)) xor (A(12) and B(116)) xor (A(13) and B(115)) xor (A(14) and B(114)) xor (A(15) and B(113)) xor (A(16) and B(112)) xor (A(17) and B(111)) xor (A(18) and B(110)) xor (A(19) and B(109)) xor (A(20) and B(108)) xor (A(21) and B(107)) xor (A(23) and B(106)) xor (A(23) and B(105)) xor (A(24) and B(104)) xor (A(25) and B(103)) xor (A(26) and B(102)) xor (A(27) and B(101)) xor (A(28) and B(100)) xor (A(29) and B(99)) xor (A(30) and B(98)) xor (A(31) and B(97)) xor (A(32) and B(96)) xor (A(33) and B(95)) xor (A(34) and B(94)) xor (A(35) and B(93)) xor (A(36) and B(92)) xor (A(37) and B(91)) xor (A(38) and B(90)) xor (A(39) and B(89)) xor (A(40) and B(88)) xor (A(41) and B(87)) xor (A(42) and B(86)) xor (A(43) and B(85)) xor (A(44) and B(84)) xor (A(45) and B(83)) xor (A(46) and B(82)) xor (A(47) and B(81)) xor (A(48) and B(80)) xor (A(49) and B(79)) xor (A(50) and B(78)) xor (A(51) and B(77)) xor (A(52) and B(76)) xor (A(53) and B(75)) xor (A(54) and B(74)) xor (A(55) and B(73)) xor (A(56) and B(72)) xor (A(57) and B(71)) xor (A(58) and B(70)) xor (A(59) and B(69)) xor (A(60) and B(68)) xor (A(61) and B(67)) xor (A(62) and B(66)) xor (A(63) and B(65)) xor (A(64) and B(64)) xor (A(65) and B(63)) xor (A(66) and B(62)) xor (A(67) and B(61)) xor (A(68) and B(60)) xor (A(69) and B(59)) xor (A(70) and B(58)) xor (A(71) and B(57)) xor (A(72) and B(56)) xor (A(73) and B(55)) xor (A(74) and B(54)) xor (A(75) and B(53)) xor (A(76) and B(52)) xor (A(77) and B(51)) xor (A(78) and B(50)) xor (A(79) and B(49)) xor (A(80) and B(48)) xor (A(81) and B(47)) xor (A(82) and B(46)) xor (A(83) and B(45)) xor (A(84) and B(44)) xor (A(85) and B(43)) xor (A(86) and B(42)) xor (A(87) and B(41)) xor (A(88) and B(40)) xor (A(89) and B(39)) xor (A(90) and B(38)) xor (A(91) and B(37)) xor (A(92) and B(36)) xor (A(93) and B(35)) xor (A(94) and B(34)) xor (A(95) and B(33)) xor (A(96) and B(32)) xor (A(97) and B(31)) xor (A(98) and B(30)) xor (A(99) and B(29)) xor (A(100) and B(28)) xor (A(101) and B(27)) xor (A(102) and B(26)) xor (A(103) and B(25)) xor (A(104) and B(24)) xor (A(105) and B(23)) xor (A(106) and B(23)) xor (A(107) and B(21)) xor (A(108) and B(20)) xor (A(109) and B(19)) xor (A(110) and B(18)) xor (A(111) and B(17)) xor (A(112) and B(16)) xor (A(113) and B(15)) xor (A(114) and B(14)) xor (A(115) and B(13)) xor (A(116) and B(12)) xor (A(117) and B(11)) xor (A(118) and B(10)) xor (A(119) and B(9)) xor (A(120) and B(8)) xor (A(121) and B(7)) xor (A(122) and B(6)) xor (A(123) and B(5)) xor (A(124) and B(4)) xor (A(125) and B(3)) xor (A(126) and B(2)) xor (A(2) and B(127)) xor (A(3) and B(126)) xor (A(4) and B(125)) xor (A(5) and B(124)) xor (A(6) and B(123)) xor (A(7) and B(122)) xor (A(8) and B(121)) xor (A(9) and B(120)) xor (A(10) and B(119)) xor (A(11) and B(118)) xor (A(12) and B(117)) xor (A(13) and B(116)) xor (A(14) and B(115)) xor (A(15) and B(114)) xor (A(16) and B(113)) xor (A(17) and B(112)) xor (A(18) and B(111)) xor (A(19) and B(110)) xor (A(20) and B(109)) xor (A(21) and B(108)) xor (A(23) and B(107)) xor (A(23) and B(106)) xor (A(24) and B(105)) xor (A(25) and B(104)) xor (A(26) and B(103)) xor (A(27) and B(102)) xor (A(28) and B(101)) xor (A(29) and B(100)) xor (A(30) and B(99)) xor (A(31) and B(98)) xor (A(32) and B(97)) xor (A(33) and B(96)) xor (A(34) and B(95)) xor (A(35) and B(94)) xor (A(36) and B(93)) xor (A(37) and B(92)) xor (A(38) and B(91)) xor (A(39) and B(90)) xor (A(40) and B(89)) xor (A(41) and B(88)) xor (A(42) and B(87)) xor (A(43) and B(86)) xor (A(44) and B(85)) xor (A(45) and B(84)) xor (A(46) and B(83)) xor (A(47) and B(82)) xor (A(48) and B(81)) xor (A(49) and B(80)) xor (A(50) and B(79)) xor (A(51) and B(78)) xor (A(52) and B(77)) xor (A(53) and B(76)) xor (A(54) and B(75)) xor (A(55) and B(74)) xor (A(56) and B(73)) xor (A(57) and B(72)) xor (A(58) and B(71)) xor (A(59) and B(70)) xor (A(60) and B(69)) xor (A(61) and B(68)) xor (A(62) and B(67)) xor (A(63) and B(66)) xor (A(64) and B(65)) xor (A(65) and B(64)) xor (A(66) and B(63)) xor (A(67) and B(62)) xor (A(68) and B(61)) xor (A(69) and B(60)) xor (A(70) and B(59)) xor (A(71) and B(58)) xor (A(72) and B(57)) xor (A(73) and B(56)) xor (A(74) and B(55)) xor (A(75) and B(54)) xor (A(76) and B(53)) xor (A(77) and B(52)) xor (A(78) and B(51)) xor (A(79) and B(50)) xor (A(80) and B(49)) xor (A(81) and B(48)) xor (A(82) and B(47)) xor (A(83) and B(46)) xor (A(84) and B(45)) xor (A(85) and B(44)) xor (A(86) and B(43)) xor (A(87) and B(42)) xor (A(88) and B(41)) xor (A(89) and B(40)) xor (A(90) and B(39)) xor (A(91) and B(38)) xor (A(92) and B(37)) xor (A(93) and B(36)) xor (A(94) and B(35)) xor (A(95) and B(34)) xor (A(96) and B(33)) xor (A(97) and B(32)) xor (A(98) and B(31)) xor (A(99) and B(30)) xor (A(100) and B(29)) xor (A(101) and B(28)) xor (A(102) and B(27)) xor (A(103) and B(26)) xor (A(104) and B(25)) xor (A(105) and B(24)) xor (A(106) and B(23)) xor (A(107) and B(23)) xor (A(108) and B(21)) xor (A(109) and B(20)) xor (A(110) and B(19)) xor (A(111) and B(18)) xor (A(112) and B(17)) xor (A(113) and B(16)) xor (A(114) and B(15)) xor (A(115) and B(14)) xor (A(116) and B(13)) xor (A(117) and B(12)) xor (A(118) and B(11)) xor (A(119) and B(10)) xor (A(120) and B(9)) xor (A(121) and B(8)) xor (A(122) and B(7)) xor (A(123) and B(6)) xor (A(124) and B(5)) xor (A(125) and B(4)) xor (A(126) and B(3)) xor (A(3) and B(127)) xor (A(4) and B(126)) xor (A(5) and B(125)) xor (A(6) and B(124)) xor (A(7) and B(123)) xor (A(8) and B(122)) xor (A(9) and B(121)) xor (A(10) and B(120)) xor (A(11) and B(119)) xor (A(12) and B(118)) xor (A(13) and B(117)) xor (A(14) and B(116)) xor (A(15) and B(115)) xor (A(16) and B(114)) xor (A(17) and B(113)) xor (A(18) and B(112)) xor (A(19) and B(111)) xor (A(20) and B(110)) xor (A(21) and B(109)) xor (A(23) and B(108)) xor (A(23) and B(107)) xor (A(24) and B(106)) xor (A(25) and B(105)) xor (A(26) and B(104)) xor (A(27) and B(103)) xor (A(28) and B(102)) xor (A(29) and B(101)) xor (A(30) and B(100)) xor (A(31) and B(99)) xor (A(32) and B(98)) xor (A(33) and B(97)) xor (A(34) and B(96)) xor (A(35) and B(95)) xor (A(36) and B(94)) xor (A(37) and B(93)) xor (A(38) and B(92)) xor (A(39) and B(91)) xor (A(40) and B(90)) xor (A(41) and B(89)) xor (A(42) and B(88)) xor (A(43) and B(87)) xor (A(44) and B(86)) xor (A(45) and B(85)) xor (A(46) and B(84)) xor (A(47) and B(83)) xor (A(48) and B(82)) xor (A(49) and B(81)) xor (A(50) and B(80)) xor (A(51) and B(79)) xor (A(52) and B(78)) xor (A(53) and B(77)) xor (A(54) and B(76)) xor (A(55) and B(75)) xor (A(56) and B(74)) xor (A(57) and B(73)) xor (A(58) and B(72)) xor (A(59) and B(71)) xor (A(60) and B(70)) xor (A(61) and B(69)) xor (A(62) and B(68)) xor (A(63) and B(67)) xor (A(64) and B(66)) xor (A(65) and B(65)) xor (A(66) and B(64)) xor (A(67) and B(63)) xor (A(68) and B(62)) xor (A(69) and B(61)) xor (A(70) and B(60)) xor (A(71) and B(59)) xor (A(72) and B(58)) xor (A(73) and B(57)) xor (A(74) and B(56)) xor (A(75) and B(55)) xor (A(76) and B(54)) xor (A(77) and B(53)) xor (A(78) and B(52)) xor (A(79) and B(51)) xor (A(80) and B(50)) xor (A(81) and B(49)) xor (A(82) and B(48)) xor (A(83) and B(47)) xor (A(84) and B(46)) xor (A(85) and B(45)) xor (A(86) and B(44)) xor (A(87) and B(43)) xor (A(88) and B(42)) xor (A(89) and B(41)) xor (A(90) and B(40)) xor (A(91) and B(39)) xor (A(92) and B(38)) xor (A(93) and B(37)) xor (A(94) and B(36)) xor (A(95) and B(35)) xor (A(96) and B(34)) xor (A(97) and B(33)) xor (A(98) and B(32)) xor (A(99) and B(31)) xor (A(100) and B(30)) xor (A(101) and B(29)) xor (A(102) and B(28)) xor (A(103) and B(27)) xor (A(104) and B(26)) xor (A(105) and B(25)) xor (A(106) and B(24)) xor (A(107) and B(23)) xor (A(108) and B(23)) xor (A(109) and B(21)) xor (A(110) and B(20)) xor (A(111) and B(19)) xor (A(112) and B(18)) xor (A(113) and B(17)) xor (A(114) and B(16)) xor (A(115) and B(15)) xor (A(116) and B(14)) xor (A(117) and B(13)) xor (A(118) and B(12)) xor (A(119) and B(11)) xor (A(120) and B(10)) xor (A(121) and B(9)) xor (A(122) and B(8)) xor (A(123) and B(7)) xor (A(124) and B(6)) xor (A(125) and B(5)) xor (A(126) and B(4)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(123)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(124)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(126));
    C(4)   <= (A(0) and B(4)) xor (A(1) and B(3)) xor (A(2) and B(2)) xor (A(3) and B(1)) xor (A(4) and B(0)) xor (A(2) and B(127)) xor (A(3) and B(126)) xor (A(4) and B(125)) xor (A(5) and B(124)) xor (A(6) and B(123)) xor (A(7) and B(122)) xor (A(8) and B(121)) xor (A(9) and B(120)) xor (A(10) and B(119)) xor (A(11) and B(118)) xor (A(12) and B(117)) xor (A(13) and B(116)) xor (A(14) and B(115)) xor (A(15) and B(114)) xor (A(16) and B(113)) xor (A(17) and B(112)) xor (A(18) and B(111)) xor (A(19) and B(110)) xor (A(20) and B(109)) xor (A(21) and B(108)) xor (A(23) and B(107)) xor (A(23) and B(106)) xor (A(24) and B(105)) xor (A(25) and B(104)) xor (A(26) and B(103)) xor (A(27) and B(102)) xor (A(28) and B(101)) xor (A(29) and B(100)) xor (A(30) and B(99)) xor (A(31) and B(98)) xor (A(32) and B(97)) xor (A(33) and B(96)) xor (A(34) and B(95)) xor (A(35) and B(94)) xor (A(36) and B(93)) xor (A(37) and B(92)) xor (A(38) and B(91)) xor (A(39) and B(90)) xor (A(40) and B(89)) xor (A(41) and B(88)) xor (A(42) and B(87)) xor (A(43) and B(86)) xor (A(44) and B(85)) xor (A(45) and B(84)) xor (A(46) and B(83)) xor (A(47) and B(82)) xor (A(48) and B(81)) xor (A(49) and B(80)) xor (A(50) and B(79)) xor (A(51) and B(78)) xor (A(52) and B(77)) xor (A(53) and B(76)) xor (A(54) and B(75)) xor (A(55) and B(74)) xor (A(56) and B(73)) xor (A(57) and B(72)) xor (A(58) and B(71)) xor (A(59) and B(70)) xor (A(60) and B(69)) xor (A(61) and B(68)) xor (A(62) and B(67)) xor (A(63) and B(66)) xor (A(64) and B(65)) xor (A(65) and B(64)) xor (A(66) and B(63)) xor (A(67) and B(62)) xor (A(68) and B(61)) xor (A(69) and B(60)) xor (A(70) and B(59)) xor (A(71) and B(58)) xor (A(72) and B(57)) xor (A(73) and B(56)) xor (A(74) and B(55)) xor (A(75) and B(54)) xor (A(76) and B(53)) xor (A(77) and B(52)) xor (A(78) and B(51)) xor (A(79) and B(50)) xor (A(80) and B(49)) xor (A(81) and B(48)) xor (A(82) and B(47)) xor (A(83) and B(46)) xor (A(84) and B(45)) xor (A(85) and B(44)) xor (A(86) and B(43)) xor (A(87) and B(42)) xor (A(88) and B(41)) xor (A(89) and B(40)) xor (A(90) and B(39)) xor (A(91) and B(38)) xor (A(92) and B(37)) xor (A(93) and B(36)) xor (A(94) and B(35)) xor (A(95) and B(34)) xor (A(96) and B(33)) xor (A(97) and B(32)) xor (A(98) and B(31)) xor (A(99) and B(30)) xor (A(100) and B(29)) xor (A(101) and B(28)) xor (A(102) and B(27)) xor (A(103) and B(26)) xor (A(104) and B(25)) xor (A(105) and B(24)) xor (A(106) and B(23)) xor (A(107) and B(23)) xor (A(108) and B(21)) xor (A(109) and B(20)) xor (A(110) and B(19)) xor (A(111) and B(18)) xor (A(112) and B(17)) xor (A(113) and B(16)) xor (A(114) and B(15)) xor (A(115) and B(14)) xor (A(116) and B(13)) xor (A(117) and B(12)) xor (A(118) and B(11)) xor (A(119) and B(10)) xor (A(120) and B(9)) xor (A(121) and B(8)) xor (A(122) and B(7)) xor (A(123) and B(6)) xor (A(124) and B(5)) xor (A(125) and B(4)) xor (A(126) and B(3)) xor (A(3) and B(127)) xor (A(4) and B(126)) xor (A(5) and B(125)) xor (A(6) and B(124)) xor (A(7) and B(123)) xor (A(8) and B(122)) xor (A(9) and B(121)) xor (A(10) and B(120)) xor (A(11) and B(119)) xor (A(12) and B(118)) xor (A(13) and B(117)) xor (A(14) and B(116)) xor (A(15) and B(115)) xor (A(16) and B(114)) xor (A(17) and B(113)) xor (A(18) and B(112)) xor (A(19) and B(111)) xor (A(20) and B(110)) xor (A(21) and B(109)) xor (A(23) and B(108)) xor (A(23) and B(107)) xor (A(24) and B(106)) xor (A(25) and B(105)) xor (A(26) and B(104)) xor (A(27) and B(103)) xor (A(28) and B(102)) xor (A(29) and B(101)) xor (A(30) and B(100)) xor (A(31) and B(99)) xor (A(32) and B(98)) xor (A(33) and B(97)) xor (A(34) and B(96)) xor (A(35) and B(95)) xor (A(36) and B(94)) xor (A(37) and B(93)) xor (A(38) and B(92)) xor (A(39) and B(91)) xor (A(40) and B(90)) xor (A(41) and B(89)) xor (A(42) and B(88)) xor (A(43) and B(87)) xor (A(44) and B(86)) xor (A(45) and B(85)) xor (A(46) and B(84)) xor (A(47) and B(83)) xor (A(48) and B(82)) xor (A(49) and B(81)) xor (A(50) and B(80)) xor (A(51) and B(79)) xor (A(52) and B(78)) xor (A(53) and B(77)) xor (A(54) and B(76)) xor (A(55) and B(75)) xor (A(56) and B(74)) xor (A(57) and B(73)) xor (A(58) and B(72)) xor (A(59) and B(71)) xor (A(60) and B(70)) xor (A(61) and B(69)) xor (A(62) and B(68)) xor (A(63) and B(67)) xor (A(64) and B(66)) xor (A(65) and B(65)) xor (A(66) and B(64)) xor (A(67) and B(63)) xor (A(68) and B(62)) xor (A(69) and B(61)) xor (A(70) and B(60)) xor (A(71) and B(59)) xor (A(72) and B(58)) xor (A(73) and B(57)) xor (A(74) and B(56)) xor (A(75) and B(55)) xor (A(76) and B(54)) xor (A(77) and B(53)) xor (A(78) and B(52)) xor (A(79) and B(51)) xor (A(80) and B(50)) xor (A(81) and B(49)) xor (A(82) and B(48)) xor (A(83) and B(47)) xor (A(84) and B(46)) xor (A(85) and B(45)) xor (A(86) and B(44)) xor (A(87) and B(43)) xor (A(88) and B(42)) xor (A(89) and B(41)) xor (A(90) and B(40)) xor (A(91) and B(39)) xor (A(92) and B(38)) xor (A(93) and B(37)) xor (A(94) and B(36)) xor (A(95) and B(35)) xor (A(96) and B(34)) xor (A(97) and B(33)) xor (A(98) and B(32)) xor (A(99) and B(31)) xor (A(100) and B(30)) xor (A(101) and B(29)) xor (A(102) and B(28)) xor (A(103) and B(27)) xor (A(104) and B(26)) xor (A(105) and B(25)) xor (A(106) and B(24)) xor (A(107) and B(23)) xor (A(108) and B(23)) xor (A(109) and B(21)) xor (A(110) and B(20)) xor (A(111) and B(19)) xor (A(112) and B(18)) xor (A(113) and B(17)) xor (A(114) and B(16)) xor (A(115) and B(15)) xor (A(116) and B(14)) xor (A(117) and B(13)) xor (A(118) and B(12)) xor (A(119) and B(11)) xor (A(120) and B(10)) xor (A(121) and B(9)) xor (A(122) and B(8)) xor (A(123) and B(7)) xor (A(124) and B(6)) xor (A(125) and B(5)) xor (A(126) and B(4)) xor (A(4) and B(127)) xor (A(5) and B(126)) xor (A(6) and B(125)) xor (A(7) and B(124)) xor (A(8) and B(123)) xor (A(9) and B(122)) xor (A(10) and B(121)) xor (A(11) and B(120)) xor (A(12) and B(119)) xor (A(13) and B(118)) xor (A(14) and B(117)) xor (A(15) and B(116)) xor (A(16) and B(115)) xor (A(17) and B(114)) xor (A(18) and B(113)) xor (A(19) and B(112)) xor (A(20) and B(111)) xor (A(21) and B(110)) xor (A(23) and B(109)) xor (A(23) and B(108)) xor (A(24) and B(107)) xor (A(25) and B(106)) xor (A(26) and B(105)) xor (A(27) and B(104)) xor (A(28) and B(103)) xor (A(29) and B(102)) xor (A(30) and B(101)) xor (A(31) and B(100)) xor (A(32) and B(99)) xor (A(33) and B(98)) xor (A(34) and B(97)) xor (A(35) and B(96)) xor (A(36) and B(95)) xor (A(37) and B(94)) xor (A(38) and B(93)) xor (A(39) and B(92)) xor (A(40) and B(91)) xor (A(41) and B(90)) xor (A(42) and B(89)) xor (A(43) and B(88)) xor (A(44) and B(87)) xor (A(45) and B(86)) xor (A(46) and B(85)) xor (A(47) and B(84)) xor (A(48) and B(83)) xor (A(49) and B(82)) xor (A(50) and B(81)) xor (A(51) and B(80)) xor (A(52) and B(79)) xor (A(53) and B(78)) xor (A(54) and B(77)) xor (A(55) and B(76)) xor (A(56) and B(75)) xor (A(57) and B(74)) xor (A(58) and B(73)) xor (A(59) and B(72)) xor (A(60) and B(71)) xor (A(61) and B(70)) xor (A(62) and B(69)) xor (A(63) and B(68)) xor (A(64) and B(67)) xor (A(65) and B(66)) xor (A(66) and B(65)) xor (A(67) and B(64)) xor (A(68) and B(63)) xor (A(69) and B(62)) xor (A(70) and B(61)) xor (A(71) and B(60)) xor (A(72) and B(59)) xor (A(73) and B(58)) xor (A(74) and B(57)) xor (A(75) and B(56)) xor (A(76) and B(55)) xor (A(77) and B(54)) xor (A(78) and B(53)) xor (A(79) and B(52)) xor (A(80) and B(51)) xor (A(81) and B(50)) xor (A(82) and B(49)) xor (A(83) and B(48)) xor (A(84) and B(47)) xor (A(85) and B(46)) xor (A(86) and B(45)) xor (A(87) and B(44)) xor (A(88) and B(43)) xor (A(89) and B(42)) xor (A(90) and B(41)) xor (A(91) and B(40)) xor (A(92) and B(39)) xor (A(93) and B(38)) xor (A(94) and B(37)) xor (A(95) and B(36)) xor (A(96) and B(35)) xor (A(97) and B(34)) xor (A(98) and B(33)) xor (A(99) and B(32)) xor (A(100) and B(31)) xor (A(101) and B(30)) xor (A(102) and B(29)) xor (A(103) and B(28)) xor (A(104) and B(27)) xor (A(105) and B(26)) xor (A(106) and B(25)) xor (A(107) and B(24)) xor (A(108) and B(23)) xor (A(109) and B(23)) xor (A(110) and B(21)) xor (A(111) and B(20)) xor (A(112) and B(19)) xor (A(113) and B(18)) xor (A(114) and B(17)) xor (A(115) and B(16)) xor (A(116) and B(15)) xor (A(117) and B(14)) xor (A(118) and B(13)) xor (A(119) and B(12)) xor (A(120) and B(11)) xor (A(121) and B(10)) xor (A(122) and B(9)) xor (A(123) and B(8)) xor (A(124) and B(7)) xor (A(125) and B(6)) xor (A(126) and B(5)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(124)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(125)) xor (A(125) and B(127)) xor (A(126) and B(127));
    C(5)   <= (A(0) and B(5)) xor (A(1) and B(4)) xor (A(2) and B(3)) xor (A(3) and B(2)) xor (A(4) and B(1)) xor (A(5) and B(0)) xor (A(3) and B(127)) xor (A(4) and B(126)) xor (A(5) and B(125)) xor (A(6) and B(124)) xor (A(7) and B(123)) xor (A(8) and B(122)) xor (A(9) and B(121)) xor (A(10) and B(120)) xor (A(11) and B(119)) xor (A(12) and B(118)) xor (A(13) and B(117)) xor (A(14) and B(116)) xor (A(15) and B(115)) xor (A(16) and B(114)) xor (A(17) and B(113)) xor (A(18) and B(112)) xor (A(19) and B(111)) xor (A(20) and B(110)) xor (A(21) and B(109)) xor (A(23) and B(108)) xor (A(23) and B(107)) xor (A(24) and B(106)) xor (A(25) and B(105)) xor (A(26) and B(104)) xor (A(27) and B(103)) xor (A(28) and B(102)) xor (A(29) and B(101)) xor (A(30) and B(100)) xor (A(31) and B(99)) xor (A(32) and B(98)) xor (A(33) and B(97)) xor (A(34) and B(96)) xor (A(35) and B(95)) xor (A(36) and B(94)) xor (A(37) and B(93)) xor (A(38) and B(92)) xor (A(39) and B(91)) xor (A(40) and B(90)) xor (A(41) and B(89)) xor (A(42) and B(88)) xor (A(43) and B(87)) xor (A(44) and B(86)) xor (A(45) and B(85)) xor (A(46) and B(84)) xor (A(47) and B(83)) xor (A(48) and B(82)) xor (A(49) and B(81)) xor (A(50) and B(80)) xor (A(51) and B(79)) xor (A(52) and B(78)) xor (A(53) and B(77)) xor (A(54) and B(76)) xor (A(55) and B(75)) xor (A(56) and B(74)) xor (A(57) and B(73)) xor (A(58) and B(72)) xor (A(59) and B(71)) xor (A(60) and B(70)) xor (A(61) and B(69)) xor (A(62) and B(68)) xor (A(63) and B(67)) xor (A(64) and B(66)) xor (A(65) and B(65)) xor (A(66) and B(64)) xor (A(67) and B(63)) xor (A(68) and B(62)) xor (A(69) and B(61)) xor (A(70) and B(60)) xor (A(71) and B(59)) xor (A(72) and B(58)) xor (A(73) and B(57)) xor (A(74) and B(56)) xor (A(75) and B(55)) xor (A(76) and B(54)) xor (A(77) and B(53)) xor (A(78) and B(52)) xor (A(79) and B(51)) xor (A(80) and B(50)) xor (A(81) and B(49)) xor (A(82) and B(48)) xor (A(83) and B(47)) xor (A(84) and B(46)) xor (A(85) and B(45)) xor (A(86) and B(44)) xor (A(87) and B(43)) xor (A(88) and B(42)) xor (A(89) and B(41)) xor (A(90) and B(40)) xor (A(91) and B(39)) xor (A(92) and B(38)) xor (A(93) and B(37)) xor (A(94) and B(36)) xor (A(95) and B(35)) xor (A(96) and B(34)) xor (A(97) and B(33)) xor (A(98) and B(32)) xor (A(99) and B(31)) xor (A(100) and B(30)) xor (A(101) and B(29)) xor (A(102) and B(28)) xor (A(103) and B(27)) xor (A(104) and B(26)) xor (A(105) and B(25)) xor (A(106) and B(24)) xor (A(107) and B(23)) xor (A(108) and B(23)) xor (A(109) and B(21)) xor (A(110) and B(20)) xor (A(111) and B(19)) xor (A(112) and B(18)) xor (A(113) and B(17)) xor (A(114) and B(16)) xor (A(115) and B(15)) xor (A(116) and B(14)) xor (A(117) and B(13)) xor (A(118) and B(12)) xor (A(119) and B(11)) xor (A(120) and B(10)) xor (A(121) and B(9)) xor (A(122) and B(8)) xor (A(123) and B(7)) xor (A(124) and B(6)) xor (A(125) and B(5)) xor (A(126) and B(4)) xor (A(4) and B(127)) xor (A(5) and B(126)) xor (A(6) and B(125)) xor (A(7) and B(124)) xor (A(8) and B(123)) xor (A(9) and B(122)) xor (A(10) and B(121)) xor (A(11) and B(120)) xor (A(12) and B(119)) xor (A(13) and B(118)) xor (A(14) and B(117)) xor (A(15) and B(116)) xor (A(16) and B(115)) xor (A(17) and B(114)) xor (A(18) and B(113)) xor (A(19) and B(112)) xor (A(20) and B(111)) xor (A(21) and B(110)) xor (A(23) and B(109)) xor (A(23) and B(108)) xor (A(24) and B(107)) xor (A(25) and B(106)) xor (A(26) and B(105)) xor (A(27) and B(104)) xor (A(28) and B(103)) xor (A(29) and B(102)) xor (A(30) and B(101)) xor (A(31) and B(100)) xor (A(32) and B(99)) xor (A(33) and B(98)) xor (A(34) and B(97)) xor (A(35) and B(96)) xor (A(36) and B(95)) xor (A(37) and B(94)) xor (A(38) and B(93)) xor (A(39) and B(92)) xor (A(40) and B(91)) xor (A(41) and B(90)) xor (A(42) and B(89)) xor (A(43) and B(88)) xor (A(44) and B(87)) xor (A(45) and B(86)) xor (A(46) and B(85)) xor (A(47) and B(84)) xor (A(48) and B(83)) xor (A(49) and B(82)) xor (A(50) and B(81)) xor (A(51) and B(80)) xor (A(52) and B(79)) xor (A(53) and B(78)) xor (A(54) and B(77)) xor (A(55) and B(76)) xor (A(56) and B(75)) xor (A(57) and B(74)) xor (A(58) and B(73)) xor (A(59) and B(72)) xor (A(60) and B(71)) xor (A(61) and B(70)) xor (A(62) and B(69)) xor (A(63) and B(68)) xor (A(64) and B(67)) xor (A(65) and B(66)) xor (A(66) and B(65)) xor (A(67) and B(64)) xor (A(68) and B(63)) xor (A(69) and B(62)) xor (A(70) and B(61)) xor (A(71) and B(60)) xor (A(72) and B(59)) xor (A(73) and B(58)) xor (A(74) and B(57)) xor (A(75) and B(56)) xor (A(76) and B(55)) xor (A(77) and B(54)) xor (A(78) and B(53)) xor (A(79) and B(52)) xor (A(80) and B(51)) xor (A(81) and B(50)) xor (A(82) and B(49)) xor (A(83) and B(48)) xor (A(84) and B(47)) xor (A(85) and B(46)) xor (A(86) and B(45)) xor (A(87) and B(44)) xor (A(88) and B(43)) xor (A(89) and B(42)) xor (A(90) and B(41)) xor (A(91) and B(40)) xor (A(92) and B(39)) xor (A(93) and B(38)) xor (A(94) and B(37)) xor (A(95) and B(36)) xor (A(96) and B(35)) xor (A(97) and B(34)) xor (A(98) and B(33)) xor (A(99) and B(32)) xor (A(100) and B(31)) xor (A(101) and B(30)) xor (A(102) and B(29)) xor (A(103) and B(28)) xor (A(104) and B(27)) xor (A(105) and B(26)) xor (A(106) and B(25)) xor (A(107) and B(24)) xor (A(108) and B(23)) xor (A(109) and B(23)) xor (A(110) and B(21)) xor (A(111) and B(20)) xor (A(112) and B(19)) xor (A(113) and B(18)) xor (A(114) and B(17)) xor (A(115) and B(16)) xor (A(116) and B(15)) xor (A(117) and B(14)) xor (A(118) and B(13)) xor (A(119) and B(12)) xor (A(120) and B(11)) xor (A(121) and B(10)) xor (A(122) and B(9)) xor (A(123) and B(8)) xor (A(124) and B(7)) xor (A(125) and B(6)) xor (A(126) and B(5)) xor (A(5) and B(127)) xor (A(6) and B(126)) xor (A(7) and B(125)) xor (A(8) and B(124)) xor (A(9) and B(123)) xor (A(10) and B(122)) xor (A(11) and B(121)) xor (A(12) and B(120)) xor (A(13) and B(119)) xor (A(14) and B(118)) xor (A(15) and B(117)) xor (A(16) and B(116)) xor (A(17) and B(115)) xor (A(18) and B(114)) xor (A(19) and B(113)) xor (A(20) and B(112)) xor (A(21) and B(111)) xor (A(23) and B(110)) xor (A(23) and B(109)) xor (A(24) and B(108)) xor (A(25) and B(107)) xor (A(26) and B(106)) xor (A(27) and B(105)) xor (A(28) and B(104)) xor (A(29) and B(103)) xor (A(30) and B(102)) xor (A(31) and B(101)) xor (A(32) and B(100)) xor (A(33) and B(99)) xor (A(34) and B(98)) xor (A(35) and B(97)) xor (A(36) and B(96)) xor (A(37) and B(95)) xor (A(38) and B(94)) xor (A(39) and B(93)) xor (A(40) and B(92)) xor (A(41) and B(91)) xor (A(42) and B(90)) xor (A(43) and B(89)) xor (A(44) and B(88)) xor (A(45) and B(87)) xor (A(46) and B(86)) xor (A(47) and B(85)) xor (A(48) and B(84)) xor (A(49) and B(83)) xor (A(50) and B(82)) xor (A(51) and B(81)) xor (A(52) and B(80)) xor (A(53) and B(79)) xor (A(54) and B(78)) xor (A(55) and B(77)) xor (A(56) and B(76)) xor (A(57) and B(75)) xor (A(58) and B(74)) xor (A(59) and B(73)) xor (A(60) and B(72)) xor (A(61) and B(71)) xor (A(62) and B(70)) xor (A(63) and B(69)) xor (A(64) and B(68)) xor (A(65) and B(67)) xor (A(66) and B(66)) xor (A(67) and B(65)) xor (A(68) and B(64)) xor (A(69) and B(63)) xor (A(70) and B(62)) xor (A(71) and B(61)) xor (A(72) and B(60)) xor (A(73) and B(59)) xor (A(74) and B(58)) xor (A(75) and B(57)) xor (A(76) and B(56)) xor (A(77) and B(55)) xor (A(78) and B(54)) xor (A(79) and B(53)) xor (A(80) and B(52)) xor (A(81) and B(51)) xor (A(82) and B(50)) xor (A(83) and B(49)) xor (A(84) and B(48)) xor (A(85) and B(47)) xor (A(86) and B(46)) xor (A(87) and B(45)) xor (A(88) and B(44)) xor (A(89) and B(43)) xor (A(90) and B(42)) xor (A(91) and B(41)) xor (A(92) and B(40)) xor (A(93) and B(39)) xor (A(94) and B(38)) xor (A(95) and B(37)) xor (A(96) and B(36)) xor (A(97) and B(35)) xor (A(98) and B(34)) xor (A(99) and B(33)) xor (A(100) and B(32)) xor (A(101) and B(31)) xor (A(102) and B(30)) xor (A(103) and B(29)) xor (A(104) and B(28)) xor (A(105) and B(27)) xor (A(106) and B(26)) xor (A(107) and B(25)) xor (A(108) and B(24)) xor (A(109) and B(23)) xor (A(110) and B(23)) xor (A(111) and B(21)) xor (A(112) and B(20)) xor (A(113) and B(19)) xor (A(114) and B(18)) xor (A(115) and B(17)) xor (A(116) and B(16)) xor (A(117) and B(15)) xor (A(118) and B(14)) xor (A(119) and B(13)) xor (A(120) and B(12)) xor (A(121) and B(11)) xor (A(122) and B(10)) xor (A(123) and B(9)) xor (A(124) and B(8)) xor (A(125) and B(7)) xor (A(126) and B(6)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(125)) xor (A(125) and B(127)) xor (A(126) and B(126)) xor (A(126) and B(127));
    C(6)   <= (A(0) and B(6)) xor (A(1) and B(5)) xor (A(2) and B(4)) xor (A(3) and B(3)) xor (A(4) and B(2)) xor (A(5) and B(1)) xor (A(6) and B(0)) xor (A(4) and B(127)) xor (A(5) and B(126)) xor (A(6) and B(125)) xor (A(7) and B(124)) xor (A(8) and B(123)) xor (A(9) and B(122)) xor (A(10) and B(121)) xor (A(11) and B(120)) xor (A(12) and B(119)) xor (A(13) and B(118)) xor (A(14) and B(117)) xor (A(15) and B(116)) xor (A(16) and B(115)) xor (A(17) and B(114)) xor (A(18) and B(113)) xor (A(19) and B(112)) xor (A(20) and B(111)) xor (A(21) and B(110)) xor (A(23) and B(109)) xor (A(23) and B(108)) xor (A(24) and B(107)) xor (A(25) and B(106)) xor (A(26) and B(105)) xor (A(27) and B(104)) xor (A(28) and B(103)) xor (A(29) and B(102)) xor (A(30) and B(101)) xor (A(31) and B(100)) xor (A(32) and B(99)) xor (A(33) and B(98)) xor (A(34) and B(97)) xor (A(35) and B(96)) xor (A(36) and B(95)) xor (A(37) and B(94)) xor (A(38) and B(93)) xor (A(39) and B(92)) xor (A(40) and B(91)) xor (A(41) and B(90)) xor (A(42) and B(89)) xor (A(43) and B(88)) xor (A(44) and B(87)) xor (A(45) and B(86)) xor (A(46) and B(85)) xor (A(47) and B(84)) xor (A(48) and B(83)) xor (A(49) and B(82)) xor (A(50) and B(81)) xor (A(51) and B(80)) xor (A(52) and B(79)) xor (A(53) and B(78)) xor (A(54) and B(77)) xor (A(55) and B(76)) xor (A(56) and B(75)) xor (A(57) and B(74)) xor (A(58) and B(73)) xor (A(59) and B(72)) xor (A(60) and B(71)) xor (A(61) and B(70)) xor (A(62) and B(69)) xor (A(63) and B(68)) xor (A(64) and B(67)) xor (A(65) and B(66)) xor (A(66) and B(65)) xor (A(67) and B(64)) xor (A(68) and B(63)) xor (A(69) and B(62)) xor (A(70) and B(61)) xor (A(71) and B(60)) xor (A(72) and B(59)) xor (A(73) and B(58)) xor (A(74) and B(57)) xor (A(75) and B(56)) xor (A(76) and B(55)) xor (A(77) and B(54)) xor (A(78) and B(53)) xor (A(79) and B(52)) xor (A(80) and B(51)) xor (A(81) and B(50)) xor (A(82) and B(49)) xor (A(83) and B(48)) xor (A(84) and B(47)) xor (A(85) and B(46)) xor (A(86) and B(45)) xor (A(87) and B(44)) xor (A(88) and B(43)) xor (A(89) and B(42)) xor (A(90) and B(41)) xor (A(91) and B(40)) xor (A(92) and B(39)) xor (A(93) and B(38)) xor (A(94) and B(37)) xor (A(95) and B(36)) xor (A(96) and B(35)) xor (A(97) and B(34)) xor (A(98) and B(33)) xor (A(99) and B(32)) xor (A(100) and B(31)) xor (A(101) and B(30)) xor (A(102) and B(29)) xor (A(103) and B(28)) xor (A(104) and B(27)) xor (A(105) and B(26)) xor (A(106) and B(25)) xor (A(107) and B(24)) xor (A(108) and B(23)) xor (A(109) and B(23)) xor (A(110) and B(21)) xor (A(111) and B(20)) xor (A(112) and B(19)) xor (A(113) and B(18)) xor (A(114) and B(17)) xor (A(115) and B(16)) xor (A(116) and B(15)) xor (A(117) and B(14)) xor (A(118) and B(13)) xor (A(119) and B(12)) xor (A(120) and B(11)) xor (A(121) and B(10)) xor (A(122) and B(9)) xor (A(123) and B(8)) xor (A(124) and B(7)) xor (A(125) and B(6)) xor (A(126) and B(5)) xor (A(5) and B(127)) xor (A(6) and B(126)) xor (A(7) and B(125)) xor (A(8) and B(124)) xor (A(9) and B(123)) xor (A(10) and B(122)) xor (A(11) and B(121)) xor (A(12) and B(120)) xor (A(13) and B(119)) xor (A(14) and B(118)) xor (A(15) and B(117)) xor (A(16) and B(116)) xor (A(17) and B(115)) xor (A(18) and B(114)) xor (A(19) and B(113)) xor (A(20) and B(112)) xor (A(21) and B(111)) xor (A(23) and B(110)) xor (A(23) and B(109)) xor (A(24) and B(108)) xor (A(25) and B(107)) xor (A(26) and B(106)) xor (A(27) and B(105)) xor (A(28) and B(104)) xor (A(29) and B(103)) xor (A(30) and B(102)) xor (A(31) and B(101)) xor (A(32) and B(100)) xor (A(33) and B(99)) xor (A(34) and B(98)) xor (A(35) and B(97)) xor (A(36) and B(96)) xor (A(37) and B(95)) xor (A(38) and B(94)) xor (A(39) and B(93)) xor (A(40) and B(92)) xor (A(41) and B(91)) xor (A(42) and B(90)) xor (A(43) and B(89)) xor (A(44) and B(88)) xor (A(45) and B(87)) xor (A(46) and B(86)) xor (A(47) and B(85)) xor (A(48) and B(84)) xor (A(49) and B(83)) xor (A(50) and B(82)) xor (A(51) and B(81)) xor (A(52) and B(80)) xor (A(53) and B(79)) xor (A(54) and B(78)) xor (A(55) and B(77)) xor (A(56) and B(76)) xor (A(57) and B(75)) xor (A(58) and B(74)) xor (A(59) and B(73)) xor (A(60) and B(72)) xor (A(61) and B(71)) xor (A(62) and B(70)) xor (A(63) and B(69)) xor (A(64) and B(68)) xor (A(65) and B(67)) xor (A(66) and B(66)) xor (A(67) and B(65)) xor (A(68) and B(64)) xor (A(69) and B(63)) xor (A(70) and B(62)) xor (A(71) and B(61)) xor (A(72) and B(60)) xor (A(73) and B(59)) xor (A(74) and B(58)) xor (A(75) and B(57)) xor (A(76) and B(56)) xor (A(77) and B(55)) xor (A(78) and B(54)) xor (A(79) and B(53)) xor (A(80) and B(52)) xor (A(81) and B(51)) xor (A(82) and B(50)) xor (A(83) and B(49)) xor (A(84) and B(48)) xor (A(85) and B(47)) xor (A(86) and B(46)) xor (A(87) and B(45)) xor (A(88) and B(44)) xor (A(89) and B(43)) xor (A(90) and B(42)) xor (A(91) and B(41)) xor (A(92) and B(40)) xor (A(93) and B(39)) xor (A(94) and B(38)) xor (A(95) and B(37)) xor (A(96) and B(36)) xor (A(97) and B(35)) xor (A(98) and B(34)) xor (A(99) and B(33)) xor (A(100) and B(32)) xor (A(101) and B(31)) xor (A(102) and B(30)) xor (A(103) and B(29)) xor (A(104) and B(28)) xor (A(105) and B(27)) xor (A(106) and B(26)) xor (A(107) and B(25)) xor (A(108) and B(24)) xor (A(109) and B(23)) xor (A(110) and B(23)) xor (A(111) and B(21)) xor (A(112) and B(20)) xor (A(113) and B(19)) xor (A(114) and B(18)) xor (A(115) and B(17)) xor (A(116) and B(16)) xor (A(117) and B(15)) xor (A(118) and B(14)) xor (A(119) and B(13)) xor (A(120) and B(12)) xor (A(121) and B(11)) xor (A(122) and B(10)) xor (A(123) and B(9)) xor (A(124) and B(8)) xor (A(125) and B(7)) xor (A(126) and B(6)) xor (A(6) and B(127)) xor (A(7) and B(126)) xor (A(8) and B(125)) xor (A(9) and B(124)) xor (A(10) and B(123)) xor (A(11) and B(122)) xor (A(12) and B(121)) xor (A(13) and B(120)) xor (A(14) and B(119)) xor (A(15) and B(118)) xor (A(16) and B(117)) xor (A(17) and B(116)) xor (A(18) and B(115)) xor (A(19) and B(114)) xor (A(20) and B(113)) xor (A(21) and B(112)) xor (A(23) and B(111)) xor (A(23) and B(110)) xor (A(24) and B(109)) xor (A(25) and B(108)) xor (A(26) and B(107)) xor (A(27) and B(106)) xor (A(28) and B(105)) xor (A(29) and B(104)) xor (A(30) and B(103)) xor (A(31) and B(102)) xor (A(32) and B(101)) xor (A(33) and B(100)) xor (A(34) and B(99)) xor (A(35) and B(98)) xor (A(36) and B(97)) xor (A(37) and B(96)) xor (A(38) and B(95)) xor (A(39) and B(94)) xor (A(40) and B(93)) xor (A(41) and B(92)) xor (A(42) and B(91)) xor (A(43) and B(90)) xor (A(44) and B(89)) xor (A(45) and B(88)) xor (A(46) and B(87)) xor (A(47) and B(86)) xor (A(48) and B(85)) xor (A(49) and B(84)) xor (A(50) and B(83)) xor (A(51) and B(82)) xor (A(52) and B(81)) xor (A(53) and B(80)) xor (A(54) and B(79)) xor (A(55) and B(78)) xor (A(56) and B(77)) xor (A(57) and B(76)) xor (A(58) and B(75)) xor (A(59) and B(74)) xor (A(60) and B(73)) xor (A(61) and B(72)) xor (A(62) and B(71)) xor (A(63) and B(70)) xor (A(64) and B(69)) xor (A(65) and B(68)) xor (A(66) and B(67)) xor (A(67) and B(66)) xor (A(68) and B(65)) xor (A(69) and B(64)) xor (A(70) and B(63)) xor (A(71) and B(62)) xor (A(72) and B(61)) xor (A(73) and B(60)) xor (A(74) and B(59)) xor (A(75) and B(58)) xor (A(76) and B(57)) xor (A(77) and B(56)) xor (A(78) and B(55)) xor (A(79) and B(54)) xor (A(80) and B(53)) xor (A(81) and B(52)) xor (A(82) and B(51)) xor (A(83) and B(50)) xor (A(84) and B(49)) xor (A(85) and B(48)) xor (A(86) and B(47)) xor (A(87) and B(46)) xor (A(88) and B(45)) xor (A(89) and B(44)) xor (A(90) and B(43)) xor (A(91) and B(42)) xor (A(92) and B(41)) xor (A(93) and B(40)) xor (A(94) and B(39)) xor (A(95) and B(38)) xor (A(96) and B(37)) xor (A(97) and B(36)) xor (A(98) and B(35)) xor (A(99) and B(34)) xor (A(100) and B(33)) xor (A(101) and B(32)) xor (A(102) and B(31)) xor (A(103) and B(30)) xor (A(104) and B(29)) xor (A(105) and B(28)) xor (A(106) and B(27)) xor (A(107) and B(26)) xor (A(108) and B(25)) xor (A(109) and B(24)) xor (A(110) and B(23)) xor (A(111) and B(23)) xor (A(112) and B(21)) xor (A(113) and B(20)) xor (A(114) and B(19)) xor (A(115) and B(18)) xor (A(116) and B(17)) xor (A(117) and B(16)) xor (A(118) and B(15)) xor (A(119) and B(14)) xor (A(120) and B(13)) xor (A(121) and B(12)) xor (A(122) and B(11)) xor (A(123) and B(10)) xor (A(124) and B(9)) xor (A(125) and B(8)) xor (A(126) and B(7)) xor (A(125) and B(127)) xor (A(126) and B(126)) xor (A(126) and B(127));
    C(7)   <= (A(0) and B(7)) xor (A(1) and B(6)) xor (A(2) and B(5)) xor (A(3) and B(4)) xor (A(4) and B(3)) xor (A(5) and B(2)) xor (A(6) and B(1)) xor (A(7) and B(0)) xor (A(0) and B(127)) xor (A(1) and B(126)) xor (A(2) and B(125)) xor (A(3) and B(124)) xor (A(4) and B(123)) xor (A(5) and B(122)) xor (A(6) and B(121)) xor (A(7) and B(120)) xor (A(8) and B(119)) xor (A(9) and B(118)) xor (A(10) and B(117)) xor (A(11) and B(116)) xor (A(12) and B(115)) xor (A(13) and B(114)) xor (A(14) and B(113)) xor (A(15) and B(112)) xor (A(16) and B(111)) xor (A(17) and B(110)) xor (A(18) and B(109)) xor (A(19) and B(108)) xor (A(20) and B(107)) xor (A(21) and B(106)) xor (A(23) and B(105)) xor (A(23) and B(104)) xor (A(24) and B(103)) xor (A(25) and B(102)) xor (A(26) and B(101)) xor (A(27) and B(100)) xor (A(28) and B(99)) xor (A(29) and B(98)) xor (A(30) and B(97)) xor (A(31) and B(96)) xor (A(32) and B(95)) xor (A(33) and B(94)) xor (A(34) and B(93)) xor (A(35) and B(92)) xor (A(36) and B(91)) xor (A(37) and B(90)) xor (A(38) and B(89)) xor (A(39) and B(88)) xor (A(40) and B(87)) xor (A(41) and B(86)) xor (A(42) and B(85)) xor (A(43) and B(84)) xor (A(44) and B(83)) xor (A(45) and B(82)) xor (A(46) and B(81)) xor (A(47) and B(80)) xor (A(48) and B(79)) xor (A(49) and B(78)) xor (A(50) and B(77)) xor (A(51) and B(76)) xor (A(52) and B(75)) xor (A(53) and B(74)) xor (A(54) and B(73)) xor (A(55) and B(72)) xor (A(56) and B(71)) xor (A(57) and B(70)) xor (A(58) and B(69)) xor (A(59) and B(68)) xor (A(60) and B(67)) xor (A(61) and B(66)) xor (A(62) and B(65)) xor (A(63) and B(64)) xor (A(64) and B(63)) xor (A(65) and B(62)) xor (A(66) and B(61)) xor (A(67) and B(60)) xor (A(68) and B(59)) xor (A(69) and B(58)) xor (A(70) and B(57)) xor (A(71) and B(56)) xor (A(72) and B(55)) xor (A(73) and B(54)) xor (A(74) and B(53)) xor (A(75) and B(52)) xor (A(76) and B(51)) xor (A(77) and B(50)) xor (A(78) and B(49)) xor (A(79) and B(48)) xor (A(80) and B(47)) xor (A(81) and B(46)) xor (A(82) and B(45)) xor (A(83) and B(44)) xor (A(84) and B(43)) xor (A(85) and B(42)) xor (A(86) and B(41)) xor (A(87) and B(40)) xor (A(88) and B(39)) xor (A(89) and B(38)) xor (A(90) and B(37)) xor (A(91) and B(36)) xor (A(92) and B(35)) xor (A(93) and B(34)) xor (A(94) and B(33)) xor (A(95) and B(32)) xor (A(96) and B(31)) xor (A(97) and B(30)) xor (A(98) and B(29)) xor (A(99) and B(28)) xor (A(100) and B(27)) xor (A(101) and B(26)) xor (A(102) and B(25)) xor (A(103) and B(24)) xor (A(104) and B(23)) xor (A(105) and B(23)) xor (A(106) and B(21)) xor (A(107) and B(20)) xor (A(108) and B(19)) xor (A(109) and B(18)) xor (A(110) and B(17)) xor (A(111) and B(16)) xor (A(112) and B(15)) xor (A(113) and B(14)) xor (A(114) and B(13)) xor (A(115) and B(12)) xor (A(116) and B(11)) xor (A(117) and B(10)) xor (A(118) and B(9)) xor (A(119) and B(8)) xor (A(120) and B(7)) xor (A(121) and B(6)) xor (A(122) and B(5)) xor (A(123) and B(4)) xor (A(124) and B(3)) xor (A(125) and B(2)) xor (A(126) and B(1)) xor (A(5) and B(127)) xor (A(6) and B(126)) xor (A(7) and B(125)) xor (A(8) and B(124)) xor (A(9) and B(123)) xor (A(10) and B(122)) xor (A(11) and B(121)) xor (A(12) and B(120)) xor (A(13) and B(119)) xor (A(14) and B(118)) xor (A(15) and B(117)) xor (A(16) and B(116)) xor (A(17) and B(115)) xor (A(18) and B(114)) xor (A(19) and B(113)) xor (A(20) and B(112)) xor (A(21) and B(111)) xor (A(23) and B(110)) xor (A(23) and B(109)) xor (A(24) and B(108)) xor (A(25) and B(107)) xor (A(26) and B(106)) xor (A(27) and B(105)) xor (A(28) and B(104)) xor (A(29) and B(103)) xor (A(30) and B(102)) xor (A(31) and B(101)) xor (A(32) and B(100)) xor (A(33) and B(99)) xor (A(34) and B(98)) xor (A(35) and B(97)) xor (A(36) and B(96)) xor (A(37) and B(95)) xor (A(38) and B(94)) xor (A(39) and B(93)) xor (A(40) and B(92)) xor (A(41) and B(91)) xor (A(42) and B(90)) xor (A(43) and B(89)) xor (A(44) and B(88)) xor (A(45) and B(87)) xor (A(46) and B(86)) xor (A(47) and B(85)) xor (A(48) and B(84)) xor (A(49) and B(83)) xor (A(50) and B(82)) xor (A(51) and B(81)) xor (A(52) and B(80)) xor (A(53) and B(79)) xor (A(54) and B(78)) xor (A(55) and B(77)) xor (A(56) and B(76)) xor (A(57) and B(75)) xor (A(58) and B(74)) xor (A(59) and B(73)) xor (A(60) and B(72)) xor (A(61) and B(71)) xor (A(62) and B(70)) xor (A(63) and B(69)) xor (A(64) and B(68)) xor (A(65) and B(67)) xor (A(66) and B(66)) xor (A(67) and B(65)) xor (A(68) and B(64)) xor (A(69) and B(63)) xor (A(70) and B(62)) xor (A(71) and B(61)) xor (A(72) and B(60)) xor (A(73) and B(59)) xor (A(74) and B(58)) xor (A(75) and B(57)) xor (A(76) and B(56)) xor (A(77) and B(55)) xor (A(78) and B(54)) xor (A(79) and B(53)) xor (A(80) and B(52)) xor (A(81) and B(51)) xor (A(82) and B(50)) xor (A(83) and B(49)) xor (A(84) and B(48)) xor (A(85) and B(47)) xor (A(86) and B(46)) xor (A(87) and B(45)) xor (A(88) and B(44)) xor (A(89) and B(43)) xor (A(90) and B(42)) xor (A(91) and B(41)) xor (A(92) and B(40)) xor (A(93) and B(39)) xor (A(94) and B(38)) xor (A(95) and B(37)) xor (A(96) and B(36)) xor (A(97) and B(35)) xor (A(98) and B(34)) xor (A(99) and B(33)) xor (A(100) and B(32)) xor (A(101) and B(31)) xor (A(102) and B(30)) xor (A(103) and B(29)) xor (A(104) and B(28)) xor (A(105) and B(27)) xor (A(106) and B(26)) xor (A(107) and B(25)) xor (A(108) and B(24)) xor (A(109) and B(23)) xor (A(110) and B(23)) xor (A(111) and B(21)) xor (A(112) and B(20)) xor (A(113) and B(19)) xor (A(114) and B(18)) xor (A(115) and B(17)) xor (A(116) and B(16)) xor (A(117) and B(15)) xor (A(118) and B(14)) xor (A(119) and B(13)) xor (A(120) and B(12)) xor (A(121) and B(11)) xor (A(122) and B(10)) xor (A(123) and B(9)) xor (A(124) and B(8)) xor (A(125) and B(7)) xor (A(126) and B(6)) xor (A(6) and B(127)) xor (A(7) and B(126)) xor (A(8) and B(125)) xor (A(9) and B(124)) xor (A(10) and B(123)) xor (A(11) and B(122)) xor (A(12) and B(121)) xor (A(13) and B(120)) xor (A(14) and B(119)) xor (A(15) and B(118)) xor (A(16) and B(117)) xor (A(17) and B(116)) xor (A(18) and B(115)) xor (A(19) and B(114)) xor (A(20) and B(113)) xor (A(21) and B(112)) xor (A(23) and B(111)) xor (A(23) and B(110)) xor (A(24) and B(109)) xor (A(25) and B(108)) xor (A(26) and B(107)) xor (A(27) and B(106)) xor (A(28) and B(105)) xor (A(29) and B(104)) xor (A(30) and B(103)) xor (A(31) and B(102)) xor (A(32) and B(101)) xor (A(33) and B(100)) xor (A(34) and B(99)) xor (A(35) and B(98)) xor (A(36) and B(97)) xor (A(37) and B(96)) xor (A(38) and B(95)) xor (A(39) and B(94)) xor (A(40) and B(93)) xor (A(41) and B(92)) xor (A(42) and B(91)) xor (A(43) and B(90)) xor (A(44) and B(89)) xor (A(45) and B(88)) xor (A(46) and B(87)) xor (A(47) and B(86)) xor (A(48) and B(85)) xor (A(49) and B(84)) xor (A(50) and B(83)) xor (A(51) and B(82)) xor (A(52) and B(81)) xor (A(53) and B(80)) xor (A(54) and B(79)) xor (A(55) and B(78)) xor (A(56) and B(77)) xor (A(57) and B(76)) xor (A(58) and B(75)) xor (A(59) and B(74)) xor (A(60) and B(73)) xor (A(61) and B(72)) xor (A(62) and B(71)) xor (A(63) and B(70)) xor (A(64) and B(69)) xor (A(65) and B(68)) xor (A(66) and B(67)) xor (A(67) and B(66)) xor (A(68) and B(65)) xor (A(69) and B(64)) xor (A(70) and B(63)) xor (A(71) and B(62)) xor (A(72) and B(61)) xor (A(73) and B(60)) xor (A(74) and B(59)) xor (A(75) and B(58)) xor (A(76) and B(57)) xor (A(77) and B(56)) xor (A(78) and B(55)) xor (A(79) and B(54)) xor (A(80) and B(53)) xor (A(81) and B(52)) xor (A(82) and B(51)) xor (A(83) and B(50)) xor (A(84) and B(49)) xor (A(85) and B(48)) xor (A(86) and B(47)) xor (A(87) and B(46)) xor (A(88) and B(45)) xor (A(89) and B(44)) xor (A(90) and B(43)) xor (A(91) and B(42)) xor (A(92) and B(41)) xor (A(93) and B(40)) xor (A(94) and B(39)) xor (A(95) and B(38)) xor (A(96) and B(37)) xor (A(97) and B(36)) xor (A(98) and B(35)) xor (A(99) and B(34)) xor (A(100) and B(33)) xor (A(101) and B(32)) xor (A(102) and B(31)) xor (A(103) and B(30)) xor (A(104) and B(29)) xor (A(105) and B(28)) xor (A(106) and B(27)) xor (A(107) and B(26)) xor (A(108) and B(25)) xor (A(109) and B(24)) xor (A(110) and B(23)) xor (A(111) and B(23)) xor (A(112) and B(21)) xor (A(113) and B(20)) xor (A(114) and B(19)) xor (A(115) and B(18)) xor (A(116) and B(17)) xor (A(117) and B(16)) xor (A(118) and B(15)) xor (A(119) and B(14)) xor (A(120) and B(13)) xor (A(121) and B(12)) xor (A(122) and B(11)) xor (A(123) and B(10)) xor (A(124) and B(9)) xor (A(125) and B(8)) xor (A(126) and B(7)) xor (A(7) and B(127)) xor (A(8) and B(126)) xor (A(9) and B(125)) xor (A(10) and B(124)) xor (A(11) and B(123)) xor (A(12) and B(122)) xor (A(13) and B(121)) xor (A(14) and B(120)) xor (A(15) and B(119)) xor (A(16) and B(118)) xor (A(17) and B(117)) xor (A(18) and B(116)) xor (A(19) and B(115)) xor (A(20) and B(114)) xor (A(21) and B(113)) xor (A(23) and B(112)) xor (A(23) and B(111)) xor (A(24) and B(110)) xor (A(25) and B(109)) xor (A(26) and B(108)) xor (A(27) and B(107)) xor (A(28) and B(106)) xor (A(29) and B(105)) xor (A(30) and B(104)) xor (A(31) and B(103)) xor (A(32) and B(102)) xor (A(33) and B(101)) xor (A(34) and B(100)) xor (A(35) and B(99)) xor (A(36) and B(98)) xor (A(37) and B(97)) xor (A(38) and B(96)) xor (A(39) and B(95)) xor (A(40) and B(94)) xor (A(41) and B(93)) xor (A(42) and B(92)) xor (A(43) and B(91)) xor (A(44) and B(90)) xor (A(45) and B(89)) xor (A(46) and B(88)) xor (A(47) and B(87)) xor (A(48) and B(86)) xor (A(49) and B(85)) xor (A(50) and B(84)) xor (A(51) and B(83)) xor (A(52) and B(82)) xor (A(53) and B(81)) xor (A(54) and B(80)) xor (A(55) and B(79)) xor (A(56) and B(78)) xor (A(57) and B(77)) xor (A(58) and B(76)) xor (A(59) and B(75)) xor (A(60) and B(74)) xor (A(61) and B(73)) xor (A(62) and B(72)) xor (A(63) and B(71)) xor (A(64) and B(70)) xor (A(65) and B(69)) xor (A(66) and B(68)) xor (A(67) and B(67)) xor (A(68) and B(66)) xor (A(69) and B(65)) xor (A(70) and B(64)) xor (A(71) and B(63)) xor (A(72) and B(62)) xor (A(73) and B(61)) xor (A(74) and B(60)) xor (A(75) and B(59)) xor (A(76) and B(58)) xor (A(77) and B(57)) xor (A(78) and B(56)) xor (A(79) and B(55)) xor (A(80) and B(54)) xor (A(81) and B(53)) xor (A(82) and B(52)) xor (A(83) and B(51)) xor (A(84) and B(50)) xor (A(85) and B(49)) xor (A(86) and B(48)) xor (A(87) and B(47)) xor (A(88) and B(46)) xor (A(89) and B(45)) xor (A(90) and B(44)) xor (A(91) and B(43)) xor (A(92) and B(42)) xor (A(93) and B(41)) xor (A(94) and B(40)) xor (A(95) and B(39)) xor (A(96) and B(38)) xor (A(97) and B(37)) xor (A(98) and B(36)) xor (A(99) and B(35)) xor (A(100) and B(34)) xor (A(101) and B(33)) xor (A(102) and B(32)) xor (A(103) and B(31)) xor (A(104) and B(30)) xor (A(105) and B(29)) xor (A(106) and B(28)) xor (A(107) and B(27)) xor (A(108) and B(26)) xor (A(109) and B(25)) xor (A(110) and B(24)) xor (A(111) and B(23)) xor (A(112) and B(23)) xor (A(113) and B(21)) xor (A(114) and B(20)) xor (A(115) and B(19)) xor (A(116) and B(18)) xor (A(117) and B(17)) xor (A(118) and B(16)) xor (A(119) and B(15)) xor (A(120) and B(14)) xor (A(121) and B(13)) xor (A(122) and B(12)) xor (A(123) and B(11)) xor (A(124) and B(10)) xor (A(125) and B(9)) xor (A(126) and B(8)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(123));
    C(8)   <= (A(0) and B(8)) xor (A(1) and B(7)) xor (A(2) and B(6)) xor (A(3) and B(5)) xor (A(4) and B(4)) xor (A(5) and B(3)) xor (A(6) and B(2)) xor (A(7) and B(1)) xor (A(8) and B(0)) xor (A(1) and B(127)) xor (A(2) and B(126)) xor (A(3) and B(125)) xor (A(4) and B(124)) xor (A(5) and B(123)) xor (A(6) and B(122)) xor (A(7) and B(121)) xor (A(8) and B(120)) xor (A(9) and B(119)) xor (A(10) and B(118)) xor (A(11) and B(117)) xor (A(12) and B(116)) xor (A(13) and B(115)) xor (A(14) and B(114)) xor (A(15) and B(113)) xor (A(16) and B(112)) xor (A(17) and B(111)) xor (A(18) and B(110)) xor (A(19) and B(109)) xor (A(20) and B(108)) xor (A(21) and B(107)) xor (A(23) and B(106)) xor (A(23) and B(105)) xor (A(24) and B(104)) xor (A(25) and B(103)) xor (A(26) and B(102)) xor (A(27) and B(101)) xor (A(28) and B(100)) xor (A(29) and B(99)) xor (A(30) and B(98)) xor (A(31) and B(97)) xor (A(32) and B(96)) xor (A(33) and B(95)) xor (A(34) and B(94)) xor (A(35) and B(93)) xor (A(36) and B(92)) xor (A(37) and B(91)) xor (A(38) and B(90)) xor (A(39) and B(89)) xor (A(40) and B(88)) xor (A(41) and B(87)) xor (A(42) and B(86)) xor (A(43) and B(85)) xor (A(44) and B(84)) xor (A(45) and B(83)) xor (A(46) and B(82)) xor (A(47) and B(81)) xor (A(48) and B(80)) xor (A(49) and B(79)) xor (A(50) and B(78)) xor (A(51) and B(77)) xor (A(52) and B(76)) xor (A(53) and B(75)) xor (A(54) and B(74)) xor (A(55) and B(73)) xor (A(56) and B(72)) xor (A(57) and B(71)) xor (A(58) and B(70)) xor (A(59) and B(69)) xor (A(60) and B(68)) xor (A(61) and B(67)) xor (A(62) and B(66)) xor (A(63) and B(65)) xor (A(64) and B(64)) xor (A(65) and B(63)) xor (A(66) and B(62)) xor (A(67) and B(61)) xor (A(68) and B(60)) xor (A(69) and B(59)) xor (A(70) and B(58)) xor (A(71) and B(57)) xor (A(72) and B(56)) xor (A(73) and B(55)) xor (A(74) and B(54)) xor (A(75) and B(53)) xor (A(76) and B(52)) xor (A(77) and B(51)) xor (A(78) and B(50)) xor (A(79) and B(49)) xor (A(80) and B(48)) xor (A(81) and B(47)) xor (A(82) and B(46)) xor (A(83) and B(45)) xor (A(84) and B(44)) xor (A(85) and B(43)) xor (A(86) and B(42)) xor (A(87) and B(41)) xor (A(88) and B(40)) xor (A(89) and B(39)) xor (A(90) and B(38)) xor (A(91) and B(37)) xor (A(92) and B(36)) xor (A(93) and B(35)) xor (A(94) and B(34)) xor (A(95) and B(33)) xor (A(96) and B(32)) xor (A(97) and B(31)) xor (A(98) and B(30)) xor (A(99) and B(29)) xor (A(100) and B(28)) xor (A(101) and B(27)) xor (A(102) and B(26)) xor (A(103) and B(25)) xor (A(104) and B(24)) xor (A(105) and B(23)) xor (A(106) and B(23)) xor (A(107) and B(21)) xor (A(108) and B(20)) xor (A(109) and B(19)) xor (A(110) and B(18)) xor (A(111) and B(17)) xor (A(112) and B(16)) xor (A(113) and B(15)) xor (A(114) and B(14)) xor (A(115) and B(13)) xor (A(116) and B(12)) xor (A(117) and B(11)) xor (A(118) and B(10)) xor (A(119) and B(9)) xor (A(120) and B(8)) xor (A(121) and B(7)) xor (A(122) and B(6)) xor (A(123) and B(5)) xor (A(124) and B(4)) xor (A(125) and B(3)) xor (A(126) and B(2)) xor (A(6) and B(127)) xor (A(7) and B(126)) xor (A(8) and B(125)) xor (A(9) and B(124)) xor (A(10) and B(123)) xor (A(11) and B(122)) xor (A(12) and B(121)) xor (A(13) and B(120)) xor (A(14) and B(119)) xor (A(15) and B(118)) xor (A(16) and B(117)) xor (A(17) and B(116)) xor (A(18) and B(115)) xor (A(19) and B(114)) xor (A(20) and B(113)) xor (A(21) and B(112)) xor (A(23) and B(111)) xor (A(23) and B(110)) xor (A(24) and B(109)) xor (A(25) and B(108)) xor (A(26) and B(107)) xor (A(27) and B(106)) xor (A(28) and B(105)) xor (A(29) and B(104)) xor (A(30) and B(103)) xor (A(31) and B(102)) xor (A(32) and B(101)) xor (A(33) and B(100)) xor (A(34) and B(99)) xor (A(35) and B(98)) xor (A(36) and B(97)) xor (A(37) and B(96)) xor (A(38) and B(95)) xor (A(39) and B(94)) xor (A(40) and B(93)) xor (A(41) and B(92)) xor (A(42) and B(91)) xor (A(43) and B(90)) xor (A(44) and B(89)) xor (A(45) and B(88)) xor (A(46) and B(87)) xor (A(47) and B(86)) xor (A(48) and B(85)) xor (A(49) and B(84)) xor (A(50) and B(83)) xor (A(51) and B(82)) xor (A(52) and B(81)) xor (A(53) and B(80)) xor (A(54) and B(79)) xor (A(55) and B(78)) xor (A(56) and B(77)) xor (A(57) and B(76)) xor (A(58) and B(75)) xor (A(59) and B(74)) xor (A(60) and B(73)) xor (A(61) and B(72)) xor (A(62) and B(71)) xor (A(63) and B(70)) xor (A(64) and B(69)) xor (A(65) and B(68)) xor (A(66) and B(67)) xor (A(67) and B(66)) xor (A(68) and B(65)) xor (A(69) and B(64)) xor (A(70) and B(63)) xor (A(71) and B(62)) xor (A(72) and B(61)) xor (A(73) and B(60)) xor (A(74) and B(59)) xor (A(75) and B(58)) xor (A(76) and B(57)) xor (A(77) and B(56)) xor (A(78) and B(55)) xor (A(79) and B(54)) xor (A(80) and B(53)) xor (A(81) and B(52)) xor (A(82) and B(51)) xor (A(83) and B(50)) xor (A(84) and B(49)) xor (A(85) and B(48)) xor (A(86) and B(47)) xor (A(87) and B(46)) xor (A(88) and B(45)) xor (A(89) and B(44)) xor (A(90) and B(43)) xor (A(91) and B(42)) xor (A(92) and B(41)) xor (A(93) and B(40)) xor (A(94) and B(39)) xor (A(95) and B(38)) xor (A(96) and B(37)) xor (A(97) and B(36)) xor (A(98) and B(35)) xor (A(99) and B(34)) xor (A(100) and B(33)) xor (A(101) and B(32)) xor (A(102) and B(31)) xor (A(103) and B(30)) xor (A(104) and B(29)) xor (A(105) and B(28)) xor (A(106) and B(27)) xor (A(107) and B(26)) xor (A(108) and B(25)) xor (A(109) and B(24)) xor (A(110) and B(23)) xor (A(111) and B(23)) xor (A(112) and B(21)) xor (A(113) and B(20)) xor (A(114) and B(19)) xor (A(115) and B(18)) xor (A(116) and B(17)) xor (A(117) and B(16)) xor (A(118) and B(15)) xor (A(119) and B(14)) xor (A(120) and B(13)) xor (A(121) and B(12)) xor (A(122) and B(11)) xor (A(123) and B(10)) xor (A(124) and B(9)) xor (A(125) and B(8)) xor (A(126) and B(7)) xor (A(7) and B(127)) xor (A(8) and B(126)) xor (A(9) and B(125)) xor (A(10) and B(124)) xor (A(11) and B(123)) xor (A(12) and B(122)) xor (A(13) and B(121)) xor (A(14) and B(120)) xor (A(15) and B(119)) xor (A(16) and B(118)) xor (A(17) and B(117)) xor (A(18) and B(116)) xor (A(19) and B(115)) xor (A(20) and B(114)) xor (A(21) and B(113)) xor (A(23) and B(112)) xor (A(23) and B(111)) xor (A(24) and B(110)) xor (A(25) and B(109)) xor (A(26) and B(108)) xor (A(27) and B(107)) xor (A(28) and B(106)) xor (A(29) and B(105)) xor (A(30) and B(104)) xor (A(31) and B(103)) xor (A(32) and B(102)) xor (A(33) and B(101)) xor (A(34) and B(100)) xor (A(35) and B(99)) xor (A(36) and B(98)) xor (A(37) and B(97)) xor (A(38) and B(96)) xor (A(39) and B(95)) xor (A(40) and B(94)) xor (A(41) and B(93)) xor (A(42) and B(92)) xor (A(43) and B(91)) xor (A(44) and B(90)) xor (A(45) and B(89)) xor (A(46) and B(88)) xor (A(47) and B(87)) xor (A(48) and B(86)) xor (A(49) and B(85)) xor (A(50) and B(84)) xor (A(51) and B(83)) xor (A(52) and B(82)) xor (A(53) and B(81)) xor (A(54) and B(80)) xor (A(55) and B(79)) xor (A(56) and B(78)) xor (A(57) and B(77)) xor (A(58) and B(76)) xor (A(59) and B(75)) xor (A(60) and B(74)) xor (A(61) and B(73)) xor (A(62) and B(72)) xor (A(63) and B(71)) xor (A(64) and B(70)) xor (A(65) and B(69)) xor (A(66) and B(68)) xor (A(67) and B(67)) xor (A(68) and B(66)) xor (A(69) and B(65)) xor (A(70) and B(64)) xor (A(71) and B(63)) xor (A(72) and B(62)) xor (A(73) and B(61)) xor (A(74) and B(60)) xor (A(75) and B(59)) xor (A(76) and B(58)) xor (A(77) and B(57)) xor (A(78) and B(56)) xor (A(79) and B(55)) xor (A(80) and B(54)) xor (A(81) and B(53)) xor (A(82) and B(52)) xor (A(83) and B(51)) xor (A(84) and B(50)) xor (A(85) and B(49)) xor (A(86) and B(48)) xor (A(87) and B(47)) xor (A(88) and B(46)) xor (A(89) and B(45)) xor (A(90) and B(44)) xor (A(91) and B(43)) xor (A(92) and B(42)) xor (A(93) and B(41)) xor (A(94) and B(40)) xor (A(95) and B(39)) xor (A(96) and B(38)) xor (A(97) and B(37)) xor (A(98) and B(36)) xor (A(99) and B(35)) xor (A(100) and B(34)) xor (A(101) and B(33)) xor (A(102) and B(32)) xor (A(103) and B(31)) xor (A(104) and B(30)) xor (A(105) and B(29)) xor (A(106) and B(28)) xor (A(107) and B(27)) xor (A(108) and B(26)) xor (A(109) and B(25)) xor (A(110) and B(24)) xor (A(111) and B(23)) xor (A(112) and B(23)) xor (A(113) and B(21)) xor (A(114) and B(20)) xor (A(115) and B(19)) xor (A(116) and B(18)) xor (A(117) and B(17)) xor (A(118) and B(16)) xor (A(119) and B(15)) xor (A(120) and B(14)) xor (A(121) and B(13)) xor (A(122) and B(12)) xor (A(123) and B(11)) xor (A(124) and B(10)) xor (A(125) and B(9)) xor (A(126) and B(8)) xor (A(8) and B(127)) xor (A(9) and B(126)) xor (A(10) and B(125)) xor (A(11) and B(124)) xor (A(12) and B(123)) xor (A(13) and B(122)) xor (A(14) and B(121)) xor (A(15) and B(120)) xor (A(16) and B(119)) xor (A(17) and B(118)) xor (A(18) and B(117)) xor (A(19) and B(116)) xor (A(20) and B(115)) xor (A(21) and B(114)) xor (A(23) and B(113)) xor (A(23) and B(112)) xor (A(24) and B(111)) xor (A(25) and B(110)) xor (A(26) and B(109)) xor (A(27) and B(108)) xor (A(28) and B(107)) xor (A(29) and B(106)) xor (A(30) and B(105)) xor (A(31) and B(104)) xor (A(32) and B(103)) xor (A(33) and B(102)) xor (A(34) and B(101)) xor (A(35) and B(100)) xor (A(36) and B(99)) xor (A(37) and B(98)) xor (A(38) and B(97)) xor (A(39) and B(96)) xor (A(40) and B(95)) xor (A(41) and B(94)) xor (A(42) and B(93)) xor (A(43) and B(92)) xor (A(44) and B(91)) xor (A(45) and B(90)) xor (A(46) and B(89)) xor (A(47) and B(88)) xor (A(48) and B(87)) xor (A(49) and B(86)) xor (A(50) and B(85)) xor (A(51) and B(84)) xor (A(52) and B(83)) xor (A(53) and B(82)) xor (A(54) and B(81)) xor (A(55) and B(80)) xor (A(56) and B(79)) xor (A(57) and B(78)) xor (A(58) and B(77)) xor (A(59) and B(76)) xor (A(60) and B(75)) xor (A(61) and B(74)) xor (A(62) and B(73)) xor (A(63) and B(72)) xor (A(64) and B(71)) xor (A(65) and B(70)) xor (A(66) and B(69)) xor (A(67) and B(68)) xor (A(68) and B(67)) xor (A(69) and B(66)) xor (A(70) and B(65)) xor (A(71) and B(64)) xor (A(72) and B(63)) xor (A(73) and B(62)) xor (A(74) and B(61)) xor (A(75) and B(60)) xor (A(76) and B(59)) xor (A(77) and B(58)) xor (A(78) and B(57)) xor (A(79) and B(56)) xor (A(80) and B(55)) xor (A(81) and B(54)) xor (A(82) and B(53)) xor (A(83) and B(52)) xor (A(84) and B(51)) xor (A(85) and B(50)) xor (A(86) and B(49)) xor (A(87) and B(48)) xor (A(88) and B(47)) xor (A(89) and B(46)) xor (A(90) and B(45)) xor (A(91) and B(44)) xor (A(92) and B(43)) xor (A(93) and B(42)) xor (A(94) and B(41)) xor (A(95) and B(40)) xor (A(96) and B(39)) xor (A(97) and B(38)) xor (A(98) and B(37)) xor (A(99) and B(36)) xor (A(100) and B(35)) xor (A(101) and B(34)) xor (A(102) and B(33)) xor (A(103) and B(32)) xor (A(104) and B(31)) xor (A(105) and B(30)) xor (A(106) and B(29)) xor (A(107) and B(28)) xor (A(108) and B(27)) xor (A(109) and B(26)) xor (A(110) and B(25)) xor (A(111) and B(24)) xor (A(112) and B(23)) xor (A(113) and B(23)) xor (A(114) and B(21)) xor (A(115) and B(20)) xor (A(116) and B(19)) xor (A(117) and B(18)) xor (A(118) and B(17)) xor (A(119) and B(16)) xor (A(120) and B(15)) xor (A(121) and B(14)) xor (A(122) and B(13)) xor (A(123) and B(12)) xor (A(124) and B(11)) xor (A(125) and B(10)) xor (A(126) and B(9)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(124));
    C(9)   <= (A(0) and B(9)) xor (A(1) and B(8)) xor (A(2) and B(7)) xor (A(3) and B(6)) xor (A(4) and B(5)) xor (A(5) and B(4)) xor (A(6) and B(3)) xor (A(7) and B(2)) xor (A(8) and B(1)) xor (A(9) and B(0)) xor (A(2) and B(127)) xor (A(3) and B(126)) xor (A(4) and B(125)) xor (A(5) and B(124)) xor (A(6) and B(123)) xor (A(7) and B(122)) xor (A(8) and B(121)) xor (A(9) and B(120)) xor (A(10) and B(119)) xor (A(11) and B(118)) xor (A(12) and B(117)) xor (A(13) and B(116)) xor (A(14) and B(115)) xor (A(15) and B(114)) xor (A(16) and B(113)) xor (A(17) and B(112)) xor (A(18) and B(111)) xor (A(19) and B(110)) xor (A(20) and B(109)) xor (A(21) and B(108)) xor (A(23) and B(107)) xor (A(23) and B(106)) xor (A(24) and B(105)) xor (A(25) and B(104)) xor (A(26) and B(103)) xor (A(27) and B(102)) xor (A(28) and B(101)) xor (A(29) and B(100)) xor (A(30) and B(99)) xor (A(31) and B(98)) xor (A(32) and B(97)) xor (A(33) and B(96)) xor (A(34) and B(95)) xor (A(35) and B(94)) xor (A(36) and B(93)) xor (A(37) and B(92)) xor (A(38) and B(91)) xor (A(39) and B(90)) xor (A(40) and B(89)) xor (A(41) and B(88)) xor (A(42) and B(87)) xor (A(43) and B(86)) xor (A(44) and B(85)) xor (A(45) and B(84)) xor (A(46) and B(83)) xor (A(47) and B(82)) xor (A(48) and B(81)) xor (A(49) and B(80)) xor (A(50) and B(79)) xor (A(51) and B(78)) xor (A(52) and B(77)) xor (A(53) and B(76)) xor (A(54) and B(75)) xor (A(55) and B(74)) xor (A(56) and B(73)) xor (A(57) and B(72)) xor (A(58) and B(71)) xor (A(59) and B(70)) xor (A(60) and B(69)) xor (A(61) and B(68)) xor (A(62) and B(67)) xor (A(63) and B(66)) xor (A(64) and B(65)) xor (A(65) and B(64)) xor (A(66) and B(63)) xor (A(67) and B(62)) xor (A(68) and B(61)) xor (A(69) and B(60)) xor (A(70) and B(59)) xor (A(71) and B(58)) xor (A(72) and B(57)) xor (A(73) and B(56)) xor (A(74) and B(55)) xor (A(75) and B(54)) xor (A(76) and B(53)) xor (A(77) and B(52)) xor (A(78) and B(51)) xor (A(79) and B(50)) xor (A(80) and B(49)) xor (A(81) and B(48)) xor (A(82) and B(47)) xor (A(83) and B(46)) xor (A(84) and B(45)) xor (A(85) and B(44)) xor (A(86) and B(43)) xor (A(87) and B(42)) xor (A(88) and B(41)) xor (A(89) and B(40)) xor (A(90) and B(39)) xor (A(91) and B(38)) xor (A(92) and B(37)) xor (A(93) and B(36)) xor (A(94) and B(35)) xor (A(95) and B(34)) xor (A(96) and B(33)) xor (A(97) and B(32)) xor (A(98) and B(31)) xor (A(99) and B(30)) xor (A(100) and B(29)) xor (A(101) and B(28)) xor (A(102) and B(27)) xor (A(103) and B(26)) xor (A(104) and B(25)) xor (A(105) and B(24)) xor (A(106) and B(23)) xor (A(107) and B(23)) xor (A(108) and B(21)) xor (A(109) and B(20)) xor (A(110) and B(19)) xor (A(111) and B(18)) xor (A(112) and B(17)) xor (A(113) and B(16)) xor (A(114) and B(15)) xor (A(115) and B(14)) xor (A(116) and B(13)) xor (A(117) and B(12)) xor (A(118) and B(11)) xor (A(119) and B(10)) xor (A(120) and B(9)) xor (A(121) and B(8)) xor (A(122) and B(7)) xor (A(123) and B(6)) xor (A(124) and B(5)) xor (A(125) and B(4)) xor (A(126) and B(3)) xor (A(7) and B(127)) xor (A(8) and B(126)) xor (A(9) and B(125)) xor (A(10) and B(124)) xor (A(11) and B(123)) xor (A(12) and B(122)) xor (A(13) and B(121)) xor (A(14) and B(120)) xor (A(15) and B(119)) xor (A(16) and B(118)) xor (A(17) and B(117)) xor (A(18) and B(116)) xor (A(19) and B(115)) xor (A(20) and B(114)) xor (A(21) and B(113)) xor (A(23) and B(112)) xor (A(23) and B(111)) xor (A(24) and B(110)) xor (A(25) and B(109)) xor (A(26) and B(108)) xor (A(27) and B(107)) xor (A(28) and B(106)) xor (A(29) and B(105)) xor (A(30) and B(104)) xor (A(31) and B(103)) xor (A(32) and B(102)) xor (A(33) and B(101)) xor (A(34) and B(100)) xor (A(35) and B(99)) xor (A(36) and B(98)) xor (A(37) and B(97)) xor (A(38) and B(96)) xor (A(39) and B(95)) xor (A(40) and B(94)) xor (A(41) and B(93)) xor (A(42) and B(92)) xor (A(43) and B(91)) xor (A(44) and B(90)) xor (A(45) and B(89)) xor (A(46) and B(88)) xor (A(47) and B(87)) xor (A(48) and B(86)) xor (A(49) and B(85)) xor (A(50) and B(84)) xor (A(51) and B(83)) xor (A(52) and B(82)) xor (A(53) and B(81)) xor (A(54) and B(80)) xor (A(55) and B(79)) xor (A(56) and B(78)) xor (A(57) and B(77)) xor (A(58) and B(76)) xor (A(59) and B(75)) xor (A(60) and B(74)) xor (A(61) and B(73)) xor (A(62) and B(72)) xor (A(63) and B(71)) xor (A(64) and B(70)) xor (A(65) and B(69)) xor (A(66) and B(68)) xor (A(67) and B(67)) xor (A(68) and B(66)) xor (A(69) and B(65)) xor (A(70) and B(64)) xor (A(71) and B(63)) xor (A(72) and B(62)) xor (A(73) and B(61)) xor (A(74) and B(60)) xor (A(75) and B(59)) xor (A(76) and B(58)) xor (A(77) and B(57)) xor (A(78) and B(56)) xor (A(79) and B(55)) xor (A(80) and B(54)) xor (A(81) and B(53)) xor (A(82) and B(52)) xor (A(83) and B(51)) xor (A(84) and B(50)) xor (A(85) and B(49)) xor (A(86) and B(48)) xor (A(87) and B(47)) xor (A(88) and B(46)) xor (A(89) and B(45)) xor (A(90) and B(44)) xor (A(91) and B(43)) xor (A(92) and B(42)) xor (A(93) and B(41)) xor (A(94) and B(40)) xor (A(95) and B(39)) xor (A(96) and B(38)) xor (A(97) and B(37)) xor (A(98) and B(36)) xor (A(99) and B(35)) xor (A(100) and B(34)) xor (A(101) and B(33)) xor (A(102) and B(32)) xor (A(103) and B(31)) xor (A(104) and B(30)) xor (A(105) and B(29)) xor (A(106) and B(28)) xor (A(107) and B(27)) xor (A(108) and B(26)) xor (A(109) and B(25)) xor (A(110) and B(24)) xor (A(111) and B(23)) xor (A(112) and B(23)) xor (A(113) and B(21)) xor (A(114) and B(20)) xor (A(115) and B(19)) xor (A(116) and B(18)) xor (A(117) and B(17)) xor (A(118) and B(16)) xor (A(119) and B(15)) xor (A(120) and B(14)) xor (A(121) and B(13)) xor (A(122) and B(12)) xor (A(123) and B(11)) xor (A(124) and B(10)) xor (A(125) and B(9)) xor (A(126) and B(8)) xor (A(8) and B(127)) xor (A(9) and B(126)) xor (A(10) and B(125)) xor (A(11) and B(124)) xor (A(12) and B(123)) xor (A(13) and B(122)) xor (A(14) and B(121)) xor (A(15) and B(120)) xor (A(16) and B(119)) xor (A(17) and B(118)) xor (A(18) and B(117)) xor (A(19) and B(116)) xor (A(20) and B(115)) xor (A(21) and B(114)) xor (A(23) and B(113)) xor (A(23) and B(112)) xor (A(24) and B(111)) xor (A(25) and B(110)) xor (A(26) and B(109)) xor (A(27) and B(108)) xor (A(28) and B(107)) xor (A(29) and B(106)) xor (A(30) and B(105)) xor (A(31) and B(104)) xor (A(32) and B(103)) xor (A(33) and B(102)) xor (A(34) and B(101)) xor (A(35) and B(100)) xor (A(36) and B(99)) xor (A(37) and B(98)) xor (A(38) and B(97)) xor (A(39) and B(96)) xor (A(40) and B(95)) xor (A(41) and B(94)) xor (A(42) and B(93)) xor (A(43) and B(92)) xor (A(44) and B(91)) xor (A(45) and B(90)) xor (A(46) and B(89)) xor (A(47) and B(88)) xor (A(48) and B(87)) xor (A(49) and B(86)) xor (A(50) and B(85)) xor (A(51) and B(84)) xor (A(52) and B(83)) xor (A(53) and B(82)) xor (A(54) and B(81)) xor (A(55) and B(80)) xor (A(56) and B(79)) xor (A(57) and B(78)) xor (A(58) and B(77)) xor (A(59) and B(76)) xor (A(60) and B(75)) xor (A(61) and B(74)) xor (A(62) and B(73)) xor (A(63) and B(72)) xor (A(64) and B(71)) xor (A(65) and B(70)) xor (A(66) and B(69)) xor (A(67) and B(68)) xor (A(68) and B(67)) xor (A(69) and B(66)) xor (A(70) and B(65)) xor (A(71) and B(64)) xor (A(72) and B(63)) xor (A(73) and B(62)) xor (A(74) and B(61)) xor (A(75) and B(60)) xor (A(76) and B(59)) xor (A(77) and B(58)) xor (A(78) and B(57)) xor (A(79) and B(56)) xor (A(80) and B(55)) xor (A(81) and B(54)) xor (A(82) and B(53)) xor (A(83) and B(52)) xor (A(84) and B(51)) xor (A(85) and B(50)) xor (A(86) and B(49)) xor (A(87) and B(48)) xor (A(88) and B(47)) xor (A(89) and B(46)) xor (A(90) and B(45)) xor (A(91) and B(44)) xor (A(92) and B(43)) xor (A(93) and B(42)) xor (A(94) and B(41)) xor (A(95) and B(40)) xor (A(96) and B(39)) xor (A(97) and B(38)) xor (A(98) and B(37)) xor (A(99) and B(36)) xor (A(100) and B(35)) xor (A(101) and B(34)) xor (A(102) and B(33)) xor (A(103) and B(32)) xor (A(104) and B(31)) xor (A(105) and B(30)) xor (A(106) and B(29)) xor (A(107) and B(28)) xor (A(108) and B(27)) xor (A(109) and B(26)) xor (A(110) and B(25)) xor (A(111) and B(24)) xor (A(112) and B(23)) xor (A(113) and B(23)) xor (A(114) and B(21)) xor (A(115) and B(20)) xor (A(116) and B(19)) xor (A(117) and B(18)) xor (A(118) and B(17)) xor (A(119) and B(16)) xor (A(120) and B(15)) xor (A(121) and B(14)) xor (A(122) and B(13)) xor (A(123) and B(12)) xor (A(124) and B(11)) xor (A(125) and B(10)) xor (A(126) and B(9)) xor (A(9) and B(127)) xor (A(10) and B(126)) xor (A(11) and B(125)) xor (A(12) and B(124)) xor (A(13) and B(123)) xor (A(14) and B(122)) xor (A(15) and B(121)) xor (A(16) and B(120)) xor (A(17) and B(119)) xor (A(18) and B(118)) xor (A(19) and B(117)) xor (A(20) and B(116)) xor (A(21) and B(115)) xor (A(23) and B(114)) xor (A(23) and B(113)) xor (A(24) and B(112)) xor (A(25) and B(111)) xor (A(26) and B(110)) xor (A(27) and B(109)) xor (A(28) and B(108)) xor (A(29) and B(107)) xor (A(30) and B(106)) xor (A(31) and B(105)) xor (A(32) and B(104)) xor (A(33) and B(103)) xor (A(34) and B(102)) xor (A(35) and B(101)) xor (A(36) and B(100)) xor (A(37) and B(99)) xor (A(38) and B(98)) xor (A(39) and B(97)) xor (A(40) and B(96)) xor (A(41) and B(95)) xor (A(42) and B(94)) xor (A(43) and B(93)) xor (A(44) and B(92)) xor (A(45) and B(91)) xor (A(46) and B(90)) xor (A(47) and B(89)) xor (A(48) and B(88)) xor (A(49) and B(87)) xor (A(50) and B(86)) xor (A(51) and B(85)) xor (A(52) and B(84)) xor (A(53) and B(83)) xor (A(54) and B(82)) xor (A(55) and B(81)) xor (A(56) and B(80)) xor (A(57) and B(79)) xor (A(58) and B(78)) xor (A(59) and B(77)) xor (A(60) and B(76)) xor (A(61) and B(75)) xor (A(62) and B(74)) xor (A(63) and B(73)) xor (A(64) and B(72)) xor (A(65) and B(71)) xor (A(66) and B(70)) xor (A(67) and B(69)) xor (A(68) and B(68)) xor (A(69) and B(67)) xor (A(70) and B(66)) xor (A(71) and B(65)) xor (A(72) and B(64)) xor (A(73) and B(63)) xor (A(74) and B(62)) xor (A(75) and B(61)) xor (A(76) and B(60)) xor (A(77) and B(59)) xor (A(78) and B(58)) xor (A(79) and B(57)) xor (A(80) and B(56)) xor (A(81) and B(55)) xor (A(82) and B(54)) xor (A(83) and B(53)) xor (A(84) and B(52)) xor (A(85) and B(51)) xor (A(86) and B(50)) xor (A(87) and B(49)) xor (A(88) and B(48)) xor (A(89) and B(47)) xor (A(90) and B(46)) xor (A(91) and B(45)) xor (A(92) and B(44)) xor (A(93) and B(43)) xor (A(94) and B(42)) xor (A(95) and B(41)) xor (A(96) and B(40)) xor (A(97) and B(39)) xor (A(98) and B(38)) xor (A(99) and B(37)) xor (A(100) and B(36)) xor (A(101) and B(35)) xor (A(102) and B(34)) xor (A(103) and B(33)) xor (A(104) and B(32)) xor (A(105) and B(31)) xor (A(106) and B(30)) xor (A(107) and B(29)) xor (A(108) and B(28)) xor (A(109) and B(27)) xor (A(110) and B(26)) xor (A(111) and B(25)) xor (A(112) and B(24)) xor (A(113) and B(23)) xor (A(114) and B(23)) xor (A(115) and B(21)) xor (A(116) and B(20)) xor (A(117) and B(19)) xor (A(118) and B(18)) xor (A(119) and B(17)) xor (A(120) and B(16)) xor (A(121) and B(15)) xor (A(122) and B(14)) xor (A(123) and B(13)) xor (A(124) and B(12)) xor (A(125) and B(11)) xor (A(126) and B(10)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(125));
    C(10)  <= (A(0) and B(10)) xor (A(1) and B(9)) xor (A(2) and B(8)) xor (A(3) and B(7)) xor (A(4) and B(6)) xor (A(5) and B(5)) xor (A(6) and B(4)) xor (A(7) and B(3)) xor (A(8) and B(2)) xor (A(9) and B(1)) xor (A(10) and B(0)) xor (A(3) and B(127)) xor (A(4) and B(126)) xor (A(5) and B(125)) xor (A(6) and B(124)) xor (A(7) and B(123)) xor (A(8) and B(122)) xor (A(9) and B(121)) xor (A(10) and B(120)) xor (A(11) and B(119)) xor (A(12) and B(118)) xor (A(13) and B(117)) xor (A(14) and B(116)) xor (A(15) and B(115)) xor (A(16) and B(114)) xor (A(17) and B(113)) xor (A(18) and B(112)) xor (A(19) and B(111)) xor (A(20) and B(110)) xor (A(21) and B(109)) xor (A(23) and B(108)) xor (A(23) and B(107)) xor (A(24) and B(106)) xor (A(25) and B(105)) xor (A(26) and B(104)) xor (A(27) and B(103)) xor (A(28) and B(102)) xor (A(29) and B(101)) xor (A(30) and B(100)) xor (A(31) and B(99)) xor (A(32) and B(98)) xor (A(33) and B(97)) xor (A(34) and B(96)) xor (A(35) and B(95)) xor (A(36) and B(94)) xor (A(37) and B(93)) xor (A(38) and B(92)) xor (A(39) and B(91)) xor (A(40) and B(90)) xor (A(41) and B(89)) xor (A(42) and B(88)) xor (A(43) and B(87)) xor (A(44) and B(86)) xor (A(45) and B(85)) xor (A(46) and B(84)) xor (A(47) and B(83)) xor (A(48) and B(82)) xor (A(49) and B(81)) xor (A(50) and B(80)) xor (A(51) and B(79)) xor (A(52) and B(78)) xor (A(53) and B(77)) xor (A(54) and B(76)) xor (A(55) and B(75)) xor (A(56) and B(74)) xor (A(57) and B(73)) xor (A(58) and B(72)) xor (A(59) and B(71)) xor (A(60) and B(70)) xor (A(61) and B(69)) xor (A(62) and B(68)) xor (A(63) and B(67)) xor (A(64) and B(66)) xor (A(65) and B(65)) xor (A(66) and B(64)) xor (A(67) and B(63)) xor (A(68) and B(62)) xor (A(69) and B(61)) xor (A(70) and B(60)) xor (A(71) and B(59)) xor (A(72) and B(58)) xor (A(73) and B(57)) xor (A(74) and B(56)) xor (A(75) and B(55)) xor (A(76) and B(54)) xor (A(77) and B(53)) xor (A(78) and B(52)) xor (A(79) and B(51)) xor (A(80) and B(50)) xor (A(81) and B(49)) xor (A(82) and B(48)) xor (A(83) and B(47)) xor (A(84) and B(46)) xor (A(85) and B(45)) xor (A(86) and B(44)) xor (A(87) and B(43)) xor (A(88) and B(42)) xor (A(89) and B(41)) xor (A(90) and B(40)) xor (A(91) and B(39)) xor (A(92) and B(38)) xor (A(93) and B(37)) xor (A(94) and B(36)) xor (A(95) and B(35)) xor (A(96) and B(34)) xor (A(97) and B(33)) xor (A(98) and B(32)) xor (A(99) and B(31)) xor (A(100) and B(30)) xor (A(101) and B(29)) xor (A(102) and B(28)) xor (A(103) and B(27)) xor (A(104) and B(26)) xor (A(105) and B(25)) xor (A(106) and B(24)) xor (A(107) and B(23)) xor (A(108) and B(23)) xor (A(109) and B(21)) xor (A(110) and B(20)) xor (A(111) and B(19)) xor (A(112) and B(18)) xor (A(113) and B(17)) xor (A(114) and B(16)) xor (A(115) and B(15)) xor (A(116) and B(14)) xor (A(117) and B(13)) xor (A(118) and B(12)) xor (A(119) and B(11)) xor (A(120) and B(10)) xor (A(121) and B(9)) xor (A(122) and B(8)) xor (A(123) and B(7)) xor (A(124) and B(6)) xor (A(125) and B(5)) xor (A(126) and B(4)) xor (A(8) and B(127)) xor (A(9) and B(126)) xor (A(10) and B(125)) xor (A(11) and B(124)) xor (A(12) and B(123)) xor (A(13) and B(122)) xor (A(14) and B(121)) xor (A(15) and B(120)) xor (A(16) and B(119)) xor (A(17) and B(118)) xor (A(18) and B(117)) xor (A(19) and B(116)) xor (A(20) and B(115)) xor (A(21) and B(114)) xor (A(23) and B(113)) xor (A(23) and B(112)) xor (A(24) and B(111)) xor (A(25) and B(110)) xor (A(26) and B(109)) xor (A(27) and B(108)) xor (A(28) and B(107)) xor (A(29) and B(106)) xor (A(30) and B(105)) xor (A(31) and B(104)) xor (A(32) and B(103)) xor (A(33) and B(102)) xor (A(34) and B(101)) xor (A(35) and B(100)) xor (A(36) and B(99)) xor (A(37) and B(98)) xor (A(38) and B(97)) xor (A(39) and B(96)) xor (A(40) and B(95)) xor (A(41) and B(94)) xor (A(42) and B(93)) xor (A(43) and B(92)) xor (A(44) and B(91)) xor (A(45) and B(90)) xor (A(46) and B(89)) xor (A(47) and B(88)) xor (A(48) and B(87)) xor (A(49) and B(86)) xor (A(50) and B(85)) xor (A(51) and B(84)) xor (A(52) and B(83)) xor (A(53) and B(82)) xor (A(54) and B(81)) xor (A(55) and B(80)) xor (A(56) and B(79)) xor (A(57) and B(78)) xor (A(58) and B(77)) xor (A(59) and B(76)) xor (A(60) and B(75)) xor (A(61) and B(74)) xor (A(62) and B(73)) xor (A(63) and B(72)) xor (A(64) and B(71)) xor (A(65) and B(70)) xor (A(66) and B(69)) xor (A(67) and B(68)) xor (A(68) and B(67)) xor (A(69) and B(66)) xor (A(70) and B(65)) xor (A(71) and B(64)) xor (A(72) and B(63)) xor (A(73) and B(62)) xor (A(74) and B(61)) xor (A(75) and B(60)) xor (A(76) and B(59)) xor (A(77) and B(58)) xor (A(78) and B(57)) xor (A(79) and B(56)) xor (A(80) and B(55)) xor (A(81) and B(54)) xor (A(82) and B(53)) xor (A(83) and B(52)) xor (A(84) and B(51)) xor (A(85) and B(50)) xor (A(86) and B(49)) xor (A(87) and B(48)) xor (A(88) and B(47)) xor (A(89) and B(46)) xor (A(90) and B(45)) xor (A(91) and B(44)) xor (A(92) and B(43)) xor (A(93) and B(42)) xor (A(94) and B(41)) xor (A(95) and B(40)) xor (A(96) and B(39)) xor (A(97) and B(38)) xor (A(98) and B(37)) xor (A(99) and B(36)) xor (A(100) and B(35)) xor (A(101) and B(34)) xor (A(102) and B(33)) xor (A(103) and B(32)) xor (A(104) and B(31)) xor (A(105) and B(30)) xor (A(106) and B(29)) xor (A(107) and B(28)) xor (A(108) and B(27)) xor (A(109) and B(26)) xor (A(110) and B(25)) xor (A(111) and B(24)) xor (A(112) and B(23)) xor (A(113) and B(23)) xor (A(114) and B(21)) xor (A(115) and B(20)) xor (A(116) and B(19)) xor (A(117) and B(18)) xor (A(118) and B(17)) xor (A(119) and B(16)) xor (A(120) and B(15)) xor (A(121) and B(14)) xor (A(122) and B(13)) xor (A(123) and B(12)) xor (A(124) and B(11)) xor (A(125) and B(10)) xor (A(126) and B(9)) xor (A(9) and B(127)) xor (A(10) and B(126)) xor (A(11) and B(125)) xor (A(12) and B(124)) xor (A(13) and B(123)) xor (A(14) and B(122)) xor (A(15) and B(121)) xor (A(16) and B(120)) xor (A(17) and B(119)) xor (A(18) and B(118)) xor (A(19) and B(117)) xor (A(20) and B(116)) xor (A(21) and B(115)) xor (A(23) and B(114)) xor (A(23) and B(113)) xor (A(24) and B(112)) xor (A(25) and B(111)) xor (A(26) and B(110)) xor (A(27) and B(109)) xor (A(28) and B(108)) xor (A(29) and B(107)) xor (A(30) and B(106)) xor (A(31) and B(105)) xor (A(32) and B(104)) xor (A(33) and B(103)) xor (A(34) and B(102)) xor (A(35) and B(101)) xor (A(36) and B(100)) xor (A(37) and B(99)) xor (A(38) and B(98)) xor (A(39) and B(97)) xor (A(40) and B(96)) xor (A(41) and B(95)) xor (A(42) and B(94)) xor (A(43) and B(93)) xor (A(44) and B(92)) xor (A(45) and B(91)) xor (A(46) and B(90)) xor (A(47) and B(89)) xor (A(48) and B(88)) xor (A(49) and B(87)) xor (A(50) and B(86)) xor (A(51) and B(85)) xor (A(52) and B(84)) xor (A(53) and B(83)) xor (A(54) and B(82)) xor (A(55) and B(81)) xor (A(56) and B(80)) xor (A(57) and B(79)) xor (A(58) and B(78)) xor (A(59) and B(77)) xor (A(60) and B(76)) xor (A(61) and B(75)) xor (A(62) and B(74)) xor (A(63) and B(73)) xor (A(64) and B(72)) xor (A(65) and B(71)) xor (A(66) and B(70)) xor (A(67) and B(69)) xor (A(68) and B(68)) xor (A(69) and B(67)) xor (A(70) and B(66)) xor (A(71) and B(65)) xor (A(72) and B(64)) xor (A(73) and B(63)) xor (A(74) and B(62)) xor (A(75) and B(61)) xor (A(76) and B(60)) xor (A(77) and B(59)) xor (A(78) and B(58)) xor (A(79) and B(57)) xor (A(80) and B(56)) xor (A(81) and B(55)) xor (A(82) and B(54)) xor (A(83) and B(53)) xor (A(84) and B(52)) xor (A(85) and B(51)) xor (A(86) and B(50)) xor (A(87) and B(49)) xor (A(88) and B(48)) xor (A(89) and B(47)) xor (A(90) and B(46)) xor (A(91) and B(45)) xor (A(92) and B(44)) xor (A(93) and B(43)) xor (A(94) and B(42)) xor (A(95) and B(41)) xor (A(96) and B(40)) xor (A(97) and B(39)) xor (A(98) and B(38)) xor (A(99) and B(37)) xor (A(100) and B(36)) xor (A(101) and B(35)) xor (A(102) and B(34)) xor (A(103) and B(33)) xor (A(104) and B(32)) xor (A(105) and B(31)) xor (A(106) and B(30)) xor (A(107) and B(29)) xor (A(108) and B(28)) xor (A(109) and B(27)) xor (A(110) and B(26)) xor (A(111) and B(25)) xor (A(112) and B(24)) xor (A(113) and B(23)) xor (A(114) and B(23)) xor (A(115) and B(21)) xor (A(116) and B(20)) xor (A(117) and B(19)) xor (A(118) and B(18)) xor (A(119) and B(17)) xor (A(120) and B(16)) xor (A(121) and B(15)) xor (A(122) and B(14)) xor (A(123) and B(13)) xor (A(124) and B(12)) xor (A(125) and B(11)) xor (A(126) and B(10)) xor (A(10) and B(127)) xor (A(11) and B(126)) xor (A(12) and B(125)) xor (A(13) and B(124)) xor (A(14) and B(123)) xor (A(15) and B(122)) xor (A(16) and B(121)) xor (A(17) and B(120)) xor (A(18) and B(119)) xor (A(19) and B(118)) xor (A(20) and B(117)) xor (A(21) and B(116)) xor (A(23) and B(115)) xor (A(23) and B(114)) xor (A(24) and B(113)) xor (A(25) and B(112)) xor (A(26) and B(111)) xor (A(27) and B(110)) xor (A(28) and B(109)) xor (A(29) and B(108)) xor (A(30) and B(107)) xor (A(31) and B(106)) xor (A(32) and B(105)) xor (A(33) and B(104)) xor (A(34) and B(103)) xor (A(35) and B(102)) xor (A(36) and B(101)) xor (A(37) and B(100)) xor (A(38) and B(99)) xor (A(39) and B(98)) xor (A(40) and B(97)) xor (A(41) and B(96)) xor (A(42) and B(95)) xor (A(43) and B(94)) xor (A(44) and B(93)) xor (A(45) and B(92)) xor (A(46) and B(91)) xor (A(47) and B(90)) xor (A(48) and B(89)) xor (A(49) and B(88)) xor (A(50) and B(87)) xor (A(51) and B(86)) xor (A(52) and B(85)) xor (A(53) and B(84)) xor (A(54) and B(83)) xor (A(55) and B(82)) xor (A(56) and B(81)) xor (A(57) and B(80)) xor (A(58) and B(79)) xor (A(59) and B(78)) xor (A(60) and B(77)) xor (A(61) and B(76)) xor (A(62) and B(75)) xor (A(63) and B(74)) xor (A(64) and B(73)) xor (A(65) and B(72)) xor (A(66) and B(71)) xor (A(67) and B(70)) xor (A(68) and B(69)) xor (A(69) and B(68)) xor (A(70) and B(67)) xor (A(71) and B(66)) xor (A(72) and B(65)) xor (A(73) and B(64)) xor (A(74) and B(63)) xor (A(75) and B(62)) xor (A(76) and B(61)) xor (A(77) and B(60)) xor (A(78) and B(59)) xor (A(79) and B(58)) xor (A(80) and B(57)) xor (A(81) and B(56)) xor (A(82) and B(55)) xor (A(83) and B(54)) xor (A(84) and B(53)) xor (A(85) and B(52)) xor (A(86) and B(51)) xor (A(87) and B(50)) xor (A(88) and B(49)) xor (A(89) and B(48)) xor (A(90) and B(47)) xor (A(91) and B(46)) xor (A(92) and B(45)) xor (A(93) and B(44)) xor (A(94) and B(43)) xor (A(95) and B(42)) xor (A(96) and B(41)) xor (A(97) and B(40)) xor (A(98) and B(39)) xor (A(99) and B(38)) xor (A(100) and B(37)) xor (A(101) and B(36)) xor (A(102) and B(35)) xor (A(103) and B(34)) xor (A(104) and B(33)) xor (A(105) and B(32)) xor (A(106) and B(31)) xor (A(107) and B(30)) xor (A(108) and B(29)) xor (A(109) and B(28)) xor (A(110) and B(27)) xor (A(111) and B(26)) xor (A(112) and B(25)) xor (A(113) and B(24)) xor (A(114) and B(23)) xor (A(115) and B(23)) xor (A(116) and B(21)) xor (A(117) and B(20)) xor (A(118) and B(19)) xor (A(119) and B(18)) xor (A(120) and B(17)) xor (A(121) and B(16)) xor (A(122) and B(15)) xor (A(123) and B(14)) xor (A(124) and B(13)) xor (A(125) and B(12)) xor (A(126) and B(11)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(126));
    C(11)  <= (A(0) and B(11)) xor (A(1) and B(10)) xor (A(2) and B(9)) xor (A(3) and B(8)) xor (A(4) and B(7)) xor (A(5) and B(6)) xor (A(6) and B(5)) xor (A(7) and B(4)) xor (A(8) and B(3)) xor (A(9) and B(2)) xor (A(10) and B(1)) xor (A(11) and B(0)) xor (A(4) and B(127)) xor (A(5) and B(126)) xor (A(6) and B(125)) xor (A(7) and B(124)) xor (A(8) and B(123)) xor (A(9) and B(122)) xor (A(10) and B(121)) xor (A(11) and B(120)) xor (A(12) and B(119)) xor (A(13) and B(118)) xor (A(14) and B(117)) xor (A(15) and B(116)) xor (A(16) and B(115)) xor (A(17) and B(114)) xor (A(18) and B(113)) xor (A(19) and B(112)) xor (A(20) and B(111)) xor (A(21) and B(110)) xor (A(23) and B(109)) xor (A(23) and B(108)) xor (A(24) and B(107)) xor (A(25) and B(106)) xor (A(26) and B(105)) xor (A(27) and B(104)) xor (A(28) and B(103)) xor (A(29) and B(102)) xor (A(30) and B(101)) xor (A(31) and B(100)) xor (A(32) and B(99)) xor (A(33) and B(98)) xor (A(34) and B(97)) xor (A(35) and B(96)) xor (A(36) and B(95)) xor (A(37) and B(94)) xor (A(38) and B(93)) xor (A(39) and B(92)) xor (A(40) and B(91)) xor (A(41) and B(90)) xor (A(42) and B(89)) xor (A(43) and B(88)) xor (A(44) and B(87)) xor (A(45) and B(86)) xor (A(46) and B(85)) xor (A(47) and B(84)) xor (A(48) and B(83)) xor (A(49) and B(82)) xor (A(50) and B(81)) xor (A(51) and B(80)) xor (A(52) and B(79)) xor (A(53) and B(78)) xor (A(54) and B(77)) xor (A(55) and B(76)) xor (A(56) and B(75)) xor (A(57) and B(74)) xor (A(58) and B(73)) xor (A(59) and B(72)) xor (A(60) and B(71)) xor (A(61) and B(70)) xor (A(62) and B(69)) xor (A(63) and B(68)) xor (A(64) and B(67)) xor (A(65) and B(66)) xor (A(66) and B(65)) xor (A(67) and B(64)) xor (A(68) and B(63)) xor (A(69) and B(62)) xor (A(70) and B(61)) xor (A(71) and B(60)) xor (A(72) and B(59)) xor (A(73) and B(58)) xor (A(74) and B(57)) xor (A(75) and B(56)) xor (A(76) and B(55)) xor (A(77) and B(54)) xor (A(78) and B(53)) xor (A(79) and B(52)) xor (A(80) and B(51)) xor (A(81) and B(50)) xor (A(82) and B(49)) xor (A(83) and B(48)) xor (A(84) and B(47)) xor (A(85) and B(46)) xor (A(86) and B(45)) xor (A(87) and B(44)) xor (A(88) and B(43)) xor (A(89) and B(42)) xor (A(90) and B(41)) xor (A(91) and B(40)) xor (A(92) and B(39)) xor (A(93) and B(38)) xor (A(94) and B(37)) xor (A(95) and B(36)) xor (A(96) and B(35)) xor (A(97) and B(34)) xor (A(98) and B(33)) xor (A(99) and B(32)) xor (A(100) and B(31)) xor (A(101) and B(30)) xor (A(102) and B(29)) xor (A(103) and B(28)) xor (A(104) and B(27)) xor (A(105) and B(26)) xor (A(106) and B(25)) xor (A(107) and B(24)) xor (A(108) and B(23)) xor (A(109) and B(23)) xor (A(110) and B(21)) xor (A(111) and B(20)) xor (A(112) and B(19)) xor (A(113) and B(18)) xor (A(114) and B(17)) xor (A(115) and B(16)) xor (A(116) and B(15)) xor (A(117) and B(14)) xor (A(118) and B(13)) xor (A(119) and B(12)) xor (A(120) and B(11)) xor (A(121) and B(10)) xor (A(122) and B(9)) xor (A(123) and B(8)) xor (A(124) and B(7)) xor (A(125) and B(6)) xor (A(126) and B(5)) xor (A(9) and B(127)) xor (A(10) and B(126)) xor (A(11) and B(125)) xor (A(12) and B(124)) xor (A(13) and B(123)) xor (A(14) and B(122)) xor (A(15) and B(121)) xor (A(16) and B(120)) xor (A(17) and B(119)) xor (A(18) and B(118)) xor (A(19) and B(117)) xor (A(20) and B(116)) xor (A(21) and B(115)) xor (A(23) and B(114)) xor (A(23) and B(113)) xor (A(24) and B(112)) xor (A(25) and B(111)) xor (A(26) and B(110)) xor (A(27) and B(109)) xor (A(28) and B(108)) xor (A(29) and B(107)) xor (A(30) and B(106)) xor (A(31) and B(105)) xor (A(32) and B(104)) xor (A(33) and B(103)) xor (A(34) and B(102)) xor (A(35) and B(101)) xor (A(36) and B(100)) xor (A(37) and B(99)) xor (A(38) and B(98)) xor (A(39) and B(97)) xor (A(40) and B(96)) xor (A(41) and B(95)) xor (A(42) and B(94)) xor (A(43) and B(93)) xor (A(44) and B(92)) xor (A(45) and B(91)) xor (A(46) and B(90)) xor (A(47) and B(89)) xor (A(48) and B(88)) xor (A(49) and B(87)) xor (A(50) and B(86)) xor (A(51) and B(85)) xor (A(52) and B(84)) xor (A(53) and B(83)) xor (A(54) and B(82)) xor (A(55) and B(81)) xor (A(56) and B(80)) xor (A(57) and B(79)) xor (A(58) and B(78)) xor (A(59) and B(77)) xor (A(60) and B(76)) xor (A(61) and B(75)) xor (A(62) and B(74)) xor (A(63) and B(73)) xor (A(64) and B(72)) xor (A(65) and B(71)) xor (A(66) and B(70)) xor (A(67) and B(69)) xor (A(68) and B(68)) xor (A(69) and B(67)) xor (A(70) and B(66)) xor (A(71) and B(65)) xor (A(72) and B(64)) xor (A(73) and B(63)) xor (A(74) and B(62)) xor (A(75) and B(61)) xor (A(76) and B(60)) xor (A(77) and B(59)) xor (A(78) and B(58)) xor (A(79) and B(57)) xor (A(80) and B(56)) xor (A(81) and B(55)) xor (A(82) and B(54)) xor (A(83) and B(53)) xor (A(84) and B(52)) xor (A(85) and B(51)) xor (A(86) and B(50)) xor (A(87) and B(49)) xor (A(88) and B(48)) xor (A(89) and B(47)) xor (A(90) and B(46)) xor (A(91) and B(45)) xor (A(92) and B(44)) xor (A(93) and B(43)) xor (A(94) and B(42)) xor (A(95) and B(41)) xor (A(96) and B(40)) xor (A(97) and B(39)) xor (A(98) and B(38)) xor (A(99) and B(37)) xor (A(100) and B(36)) xor (A(101) and B(35)) xor (A(102) and B(34)) xor (A(103) and B(33)) xor (A(104) and B(32)) xor (A(105) and B(31)) xor (A(106) and B(30)) xor (A(107) and B(29)) xor (A(108) and B(28)) xor (A(109) and B(27)) xor (A(110) and B(26)) xor (A(111) and B(25)) xor (A(112) and B(24)) xor (A(113) and B(23)) xor (A(114) and B(23)) xor (A(115) and B(21)) xor (A(116) and B(20)) xor (A(117) and B(19)) xor (A(118) and B(18)) xor (A(119) and B(17)) xor (A(120) and B(16)) xor (A(121) and B(15)) xor (A(122) and B(14)) xor (A(123) and B(13)) xor (A(124) and B(12)) xor (A(125) and B(11)) xor (A(126) and B(10)) xor (A(10) and B(127)) xor (A(11) and B(126)) xor (A(12) and B(125)) xor (A(13) and B(124)) xor (A(14) and B(123)) xor (A(15) and B(122)) xor (A(16) and B(121)) xor (A(17) and B(120)) xor (A(18) and B(119)) xor (A(19) and B(118)) xor (A(20) and B(117)) xor (A(21) and B(116)) xor (A(23) and B(115)) xor (A(23) and B(114)) xor (A(24) and B(113)) xor (A(25) and B(112)) xor (A(26) and B(111)) xor (A(27) and B(110)) xor (A(28) and B(109)) xor (A(29) and B(108)) xor (A(30) and B(107)) xor (A(31) and B(106)) xor (A(32) and B(105)) xor (A(33) and B(104)) xor (A(34) and B(103)) xor (A(35) and B(102)) xor (A(36) and B(101)) xor (A(37) and B(100)) xor (A(38) and B(99)) xor (A(39) and B(98)) xor (A(40) and B(97)) xor (A(41) and B(96)) xor (A(42) and B(95)) xor (A(43) and B(94)) xor (A(44) and B(93)) xor (A(45) and B(92)) xor (A(46) and B(91)) xor (A(47) and B(90)) xor (A(48) and B(89)) xor (A(49) and B(88)) xor (A(50) and B(87)) xor (A(51) and B(86)) xor (A(52) and B(85)) xor (A(53) and B(84)) xor (A(54) and B(83)) xor (A(55) and B(82)) xor (A(56) and B(81)) xor (A(57) and B(80)) xor (A(58) and B(79)) xor (A(59) and B(78)) xor (A(60) and B(77)) xor (A(61) and B(76)) xor (A(62) and B(75)) xor (A(63) and B(74)) xor (A(64) and B(73)) xor (A(65) and B(72)) xor (A(66) and B(71)) xor (A(67) and B(70)) xor (A(68) and B(69)) xor (A(69) and B(68)) xor (A(70) and B(67)) xor (A(71) and B(66)) xor (A(72) and B(65)) xor (A(73) and B(64)) xor (A(74) and B(63)) xor (A(75) and B(62)) xor (A(76) and B(61)) xor (A(77) and B(60)) xor (A(78) and B(59)) xor (A(79) and B(58)) xor (A(80) and B(57)) xor (A(81) and B(56)) xor (A(82) and B(55)) xor (A(83) and B(54)) xor (A(84) and B(53)) xor (A(85) and B(52)) xor (A(86) and B(51)) xor (A(87) and B(50)) xor (A(88) and B(49)) xor (A(89) and B(48)) xor (A(90) and B(47)) xor (A(91) and B(46)) xor (A(92) and B(45)) xor (A(93) and B(44)) xor (A(94) and B(43)) xor (A(95) and B(42)) xor (A(96) and B(41)) xor (A(97) and B(40)) xor (A(98) and B(39)) xor (A(99) and B(38)) xor (A(100) and B(37)) xor (A(101) and B(36)) xor (A(102) and B(35)) xor (A(103) and B(34)) xor (A(104) and B(33)) xor (A(105) and B(32)) xor (A(106) and B(31)) xor (A(107) and B(30)) xor (A(108) and B(29)) xor (A(109) and B(28)) xor (A(110) and B(27)) xor (A(111) and B(26)) xor (A(112) and B(25)) xor (A(113) and B(24)) xor (A(114) and B(23)) xor (A(115) and B(23)) xor (A(116) and B(21)) xor (A(117) and B(20)) xor (A(118) and B(19)) xor (A(119) and B(18)) xor (A(120) and B(17)) xor (A(121) and B(16)) xor (A(122) and B(15)) xor (A(123) and B(14)) xor (A(124) and B(13)) xor (A(125) and B(12)) xor (A(126) and B(11)) xor (A(11) and B(127)) xor (A(12) and B(126)) xor (A(13) and B(125)) xor (A(14) and B(124)) xor (A(15) and B(123)) xor (A(16) and B(122)) xor (A(17) and B(121)) xor (A(18) and B(120)) xor (A(19) and B(119)) xor (A(20) and B(118)) xor (A(21) and B(117)) xor (A(23) and B(116)) xor (A(23) and B(115)) xor (A(24) and B(114)) xor (A(25) and B(113)) xor (A(26) and B(112)) xor (A(27) and B(111)) xor (A(28) and B(110)) xor (A(29) and B(109)) xor (A(30) and B(108)) xor (A(31) and B(107)) xor (A(32) and B(106)) xor (A(33) and B(105)) xor (A(34) and B(104)) xor (A(35) and B(103)) xor (A(36) and B(102)) xor (A(37) and B(101)) xor (A(38) and B(100)) xor (A(39) and B(99)) xor (A(40) and B(98)) xor (A(41) and B(97)) xor (A(42) and B(96)) xor (A(43) and B(95)) xor (A(44) and B(94)) xor (A(45) and B(93)) xor (A(46) and B(92)) xor (A(47) and B(91)) xor (A(48) and B(90)) xor (A(49) and B(89)) xor (A(50) and B(88)) xor (A(51) and B(87)) xor (A(52) and B(86)) xor (A(53) and B(85)) xor (A(54) and B(84)) xor (A(55) and B(83)) xor (A(56) and B(82)) xor (A(57) and B(81)) xor (A(58) and B(80)) xor (A(59) and B(79)) xor (A(60) and B(78)) xor (A(61) and B(77)) xor (A(62) and B(76)) xor (A(63) and B(75)) xor (A(64) and B(74)) xor (A(65) and B(73)) xor (A(66) and B(72)) xor (A(67) and B(71)) xor (A(68) and B(70)) xor (A(69) and B(69)) xor (A(70) and B(68)) xor (A(71) and B(67)) xor (A(72) and B(66)) xor (A(73) and B(65)) xor (A(74) and B(64)) xor (A(75) and B(63)) xor (A(76) and B(62)) xor (A(77) and B(61)) xor (A(78) and B(60)) xor (A(79) and B(59)) xor (A(80) and B(58)) xor (A(81) and B(57)) xor (A(82) and B(56)) xor (A(83) and B(55)) xor (A(84) and B(54)) xor (A(85) and B(53)) xor (A(86) and B(52)) xor (A(87) and B(51)) xor (A(88) and B(50)) xor (A(89) and B(49)) xor (A(90) and B(48)) xor (A(91) and B(47)) xor (A(92) and B(46)) xor (A(93) and B(45)) xor (A(94) and B(44)) xor (A(95) and B(43)) xor (A(96) and B(42)) xor (A(97) and B(41)) xor (A(98) and B(40)) xor (A(99) and B(39)) xor (A(100) and B(38)) xor (A(101) and B(37)) xor (A(102) and B(36)) xor (A(103) and B(35)) xor (A(104) and B(34)) xor (A(105) and B(33)) xor (A(106) and B(32)) xor (A(107) and B(31)) xor (A(108) and B(30)) xor (A(109) and B(29)) xor (A(110) and B(28)) xor (A(111) and B(27)) xor (A(112) and B(26)) xor (A(113) and B(25)) xor (A(114) and B(24)) xor (A(115) and B(23)) xor (A(116) and B(23)) xor (A(117) and B(21)) xor (A(118) and B(20)) xor (A(119) and B(19)) xor (A(120) and B(18)) xor (A(121) and B(17)) xor (A(122) and B(16)) xor (A(123) and B(15)) xor (A(124) and B(14)) xor (A(125) and B(13)) xor (A(126) and B(12)) xor (A(125) and B(127)) xor (A(126) and B(127));
    C(12)  <= (A(0) and B(12)) xor (A(1) and B(11)) xor (A(2) and B(10)) xor (A(3) and B(9)) xor (A(4) and B(8)) xor (A(5) and B(7)) xor (A(6) and B(6)) xor (A(7) and B(5)) xor (A(8) and B(4)) xor (A(9) and B(3)) xor (A(10) and B(2)) xor (A(11) and B(1)) xor (A(12) and B(0)) xor (A(5) and B(127)) xor (A(6) and B(126)) xor (A(7) and B(125)) xor (A(8) and B(124)) xor (A(9) and B(123)) xor (A(10) and B(122)) xor (A(11) and B(121)) xor (A(12) and B(120)) xor (A(13) and B(119)) xor (A(14) and B(118)) xor (A(15) and B(117)) xor (A(16) and B(116)) xor (A(17) and B(115)) xor (A(18) and B(114)) xor (A(19) and B(113)) xor (A(20) and B(112)) xor (A(21) and B(111)) xor (A(23) and B(110)) xor (A(23) and B(109)) xor (A(24) and B(108)) xor (A(25) and B(107)) xor (A(26) and B(106)) xor (A(27) and B(105)) xor (A(28) and B(104)) xor (A(29) and B(103)) xor (A(30) and B(102)) xor (A(31) and B(101)) xor (A(32) and B(100)) xor (A(33) and B(99)) xor (A(34) and B(98)) xor (A(35) and B(97)) xor (A(36) and B(96)) xor (A(37) and B(95)) xor (A(38) and B(94)) xor (A(39) and B(93)) xor (A(40) and B(92)) xor (A(41) and B(91)) xor (A(42) and B(90)) xor (A(43) and B(89)) xor (A(44) and B(88)) xor (A(45) and B(87)) xor (A(46) and B(86)) xor (A(47) and B(85)) xor (A(48) and B(84)) xor (A(49) and B(83)) xor (A(50) and B(82)) xor (A(51) and B(81)) xor (A(52) and B(80)) xor (A(53) and B(79)) xor (A(54) and B(78)) xor (A(55) and B(77)) xor (A(56) and B(76)) xor (A(57) and B(75)) xor (A(58) and B(74)) xor (A(59) and B(73)) xor (A(60) and B(72)) xor (A(61) and B(71)) xor (A(62) and B(70)) xor (A(63) and B(69)) xor (A(64) and B(68)) xor (A(65) and B(67)) xor (A(66) and B(66)) xor (A(67) and B(65)) xor (A(68) and B(64)) xor (A(69) and B(63)) xor (A(70) and B(62)) xor (A(71) and B(61)) xor (A(72) and B(60)) xor (A(73) and B(59)) xor (A(74) and B(58)) xor (A(75) and B(57)) xor (A(76) and B(56)) xor (A(77) and B(55)) xor (A(78) and B(54)) xor (A(79) and B(53)) xor (A(80) and B(52)) xor (A(81) and B(51)) xor (A(82) and B(50)) xor (A(83) and B(49)) xor (A(84) and B(48)) xor (A(85) and B(47)) xor (A(86) and B(46)) xor (A(87) and B(45)) xor (A(88) and B(44)) xor (A(89) and B(43)) xor (A(90) and B(42)) xor (A(91) and B(41)) xor (A(92) and B(40)) xor (A(93) and B(39)) xor (A(94) and B(38)) xor (A(95) and B(37)) xor (A(96) and B(36)) xor (A(97) and B(35)) xor (A(98) and B(34)) xor (A(99) and B(33)) xor (A(100) and B(32)) xor (A(101) and B(31)) xor (A(102) and B(30)) xor (A(103) and B(29)) xor (A(104) and B(28)) xor (A(105) and B(27)) xor (A(106) and B(26)) xor (A(107) and B(25)) xor (A(108) and B(24)) xor (A(109) and B(23)) xor (A(110) and B(23)) xor (A(111) and B(21)) xor (A(112) and B(20)) xor (A(113) and B(19)) xor (A(114) and B(18)) xor (A(115) and B(17)) xor (A(116) and B(16)) xor (A(117) and B(15)) xor (A(118) and B(14)) xor (A(119) and B(13)) xor (A(120) and B(12)) xor (A(121) and B(11)) xor (A(122) and B(10)) xor (A(123) and B(9)) xor (A(124) and B(8)) xor (A(125) and B(7)) xor (A(126) and B(6)) xor (A(10) and B(127)) xor (A(11) and B(126)) xor (A(12) and B(125)) xor (A(13) and B(124)) xor (A(14) and B(123)) xor (A(15) and B(122)) xor (A(16) and B(121)) xor (A(17) and B(120)) xor (A(18) and B(119)) xor (A(19) and B(118)) xor (A(20) and B(117)) xor (A(21) and B(116)) xor (A(23) and B(115)) xor (A(23) and B(114)) xor (A(24) and B(113)) xor (A(25) and B(112)) xor (A(26) and B(111)) xor (A(27) and B(110)) xor (A(28) and B(109)) xor (A(29) and B(108)) xor (A(30) and B(107)) xor (A(31) and B(106)) xor (A(32) and B(105)) xor (A(33) and B(104)) xor (A(34) and B(103)) xor (A(35) and B(102)) xor (A(36) and B(101)) xor (A(37) and B(100)) xor (A(38) and B(99)) xor (A(39) and B(98)) xor (A(40) and B(97)) xor (A(41) and B(96)) xor (A(42) and B(95)) xor (A(43) and B(94)) xor (A(44) and B(93)) xor (A(45) and B(92)) xor (A(46) and B(91)) xor (A(47) and B(90)) xor (A(48) and B(89)) xor (A(49) and B(88)) xor (A(50) and B(87)) xor (A(51) and B(86)) xor (A(52) and B(85)) xor (A(53) and B(84)) xor (A(54) and B(83)) xor (A(55) and B(82)) xor (A(56) and B(81)) xor (A(57) and B(80)) xor (A(58) and B(79)) xor (A(59) and B(78)) xor (A(60) and B(77)) xor (A(61) and B(76)) xor (A(62) and B(75)) xor (A(63) and B(74)) xor (A(64) and B(73)) xor (A(65) and B(72)) xor (A(66) and B(71)) xor (A(67) and B(70)) xor (A(68) and B(69)) xor (A(69) and B(68)) xor (A(70) and B(67)) xor (A(71) and B(66)) xor (A(72) and B(65)) xor (A(73) and B(64)) xor (A(74) and B(63)) xor (A(75) and B(62)) xor (A(76) and B(61)) xor (A(77) and B(60)) xor (A(78) and B(59)) xor (A(79) and B(58)) xor (A(80) and B(57)) xor (A(81) and B(56)) xor (A(82) and B(55)) xor (A(83) and B(54)) xor (A(84) and B(53)) xor (A(85) and B(52)) xor (A(86) and B(51)) xor (A(87) and B(50)) xor (A(88) and B(49)) xor (A(89) and B(48)) xor (A(90) and B(47)) xor (A(91) and B(46)) xor (A(92) and B(45)) xor (A(93) and B(44)) xor (A(94) and B(43)) xor (A(95) and B(42)) xor (A(96) and B(41)) xor (A(97) and B(40)) xor (A(98) and B(39)) xor (A(99) and B(38)) xor (A(100) and B(37)) xor (A(101) and B(36)) xor (A(102) and B(35)) xor (A(103) and B(34)) xor (A(104) and B(33)) xor (A(105) and B(32)) xor (A(106) and B(31)) xor (A(107) and B(30)) xor (A(108) and B(29)) xor (A(109) and B(28)) xor (A(110) and B(27)) xor (A(111) and B(26)) xor (A(112) and B(25)) xor (A(113) and B(24)) xor (A(114) and B(23)) xor (A(115) and B(23)) xor (A(116) and B(21)) xor (A(117) and B(20)) xor (A(118) and B(19)) xor (A(119) and B(18)) xor (A(120) and B(17)) xor (A(121) and B(16)) xor (A(122) and B(15)) xor (A(123) and B(14)) xor (A(124) and B(13)) xor (A(125) and B(12)) xor (A(126) and B(11)) xor (A(11) and B(127)) xor (A(12) and B(126)) xor (A(13) and B(125)) xor (A(14) and B(124)) xor (A(15) and B(123)) xor (A(16) and B(122)) xor (A(17) and B(121)) xor (A(18) and B(120)) xor (A(19) and B(119)) xor (A(20) and B(118)) xor (A(21) and B(117)) xor (A(23) and B(116)) xor (A(23) and B(115)) xor (A(24) and B(114)) xor (A(25) and B(113)) xor (A(26) and B(112)) xor (A(27) and B(111)) xor (A(28) and B(110)) xor (A(29) and B(109)) xor (A(30) and B(108)) xor (A(31) and B(107)) xor (A(32) and B(106)) xor (A(33) and B(105)) xor (A(34) and B(104)) xor (A(35) and B(103)) xor (A(36) and B(102)) xor (A(37) and B(101)) xor (A(38) and B(100)) xor (A(39) and B(99)) xor (A(40) and B(98)) xor (A(41) and B(97)) xor (A(42) and B(96)) xor (A(43) and B(95)) xor (A(44) and B(94)) xor (A(45) and B(93)) xor (A(46) and B(92)) xor (A(47) and B(91)) xor (A(48) and B(90)) xor (A(49) and B(89)) xor (A(50) and B(88)) xor (A(51) and B(87)) xor (A(52) and B(86)) xor (A(53) and B(85)) xor (A(54) and B(84)) xor (A(55) and B(83)) xor (A(56) and B(82)) xor (A(57) and B(81)) xor (A(58) and B(80)) xor (A(59) and B(79)) xor (A(60) and B(78)) xor (A(61) and B(77)) xor (A(62) and B(76)) xor (A(63) and B(75)) xor (A(64) and B(74)) xor (A(65) and B(73)) xor (A(66) and B(72)) xor (A(67) and B(71)) xor (A(68) and B(70)) xor (A(69) and B(69)) xor (A(70) and B(68)) xor (A(71) and B(67)) xor (A(72) and B(66)) xor (A(73) and B(65)) xor (A(74) and B(64)) xor (A(75) and B(63)) xor (A(76) and B(62)) xor (A(77) and B(61)) xor (A(78) and B(60)) xor (A(79) and B(59)) xor (A(80) and B(58)) xor (A(81) and B(57)) xor (A(82) and B(56)) xor (A(83) and B(55)) xor (A(84) and B(54)) xor (A(85) and B(53)) xor (A(86) and B(52)) xor (A(87) and B(51)) xor (A(88) and B(50)) xor (A(89) and B(49)) xor (A(90) and B(48)) xor (A(91) and B(47)) xor (A(92) and B(46)) xor (A(93) and B(45)) xor (A(94) and B(44)) xor (A(95) and B(43)) xor (A(96) and B(42)) xor (A(97) and B(41)) xor (A(98) and B(40)) xor (A(99) and B(39)) xor (A(100) and B(38)) xor (A(101) and B(37)) xor (A(102) and B(36)) xor (A(103) and B(35)) xor (A(104) and B(34)) xor (A(105) and B(33)) xor (A(106) and B(32)) xor (A(107) and B(31)) xor (A(108) and B(30)) xor (A(109) and B(29)) xor (A(110) and B(28)) xor (A(111) and B(27)) xor (A(112) and B(26)) xor (A(113) and B(25)) xor (A(114) and B(24)) xor (A(115) and B(23)) xor (A(116) and B(23)) xor (A(117) and B(21)) xor (A(118) and B(20)) xor (A(119) and B(19)) xor (A(120) and B(18)) xor (A(121) and B(17)) xor (A(122) and B(16)) xor (A(123) and B(15)) xor (A(124) and B(14)) xor (A(125) and B(13)) xor (A(126) and B(12)) xor (A(12) and B(127)) xor (A(13) and B(126)) xor (A(14) and B(125)) xor (A(15) and B(124)) xor (A(16) and B(123)) xor (A(17) and B(122)) xor (A(18) and B(121)) xor (A(19) and B(120)) xor (A(20) and B(119)) xor (A(21) and B(118)) xor (A(23) and B(117)) xor (A(23) and B(116)) xor (A(24) and B(115)) xor (A(25) and B(114)) xor (A(26) and B(113)) xor (A(27) and B(112)) xor (A(28) and B(111)) xor (A(29) and B(110)) xor (A(30) and B(109)) xor (A(31) and B(108)) xor (A(32) and B(107)) xor (A(33) and B(106)) xor (A(34) and B(105)) xor (A(35) and B(104)) xor (A(36) and B(103)) xor (A(37) and B(102)) xor (A(38) and B(101)) xor (A(39) and B(100)) xor (A(40) and B(99)) xor (A(41) and B(98)) xor (A(42) and B(97)) xor (A(43) and B(96)) xor (A(44) and B(95)) xor (A(45) and B(94)) xor (A(46) and B(93)) xor (A(47) and B(92)) xor (A(48) and B(91)) xor (A(49) and B(90)) xor (A(50) and B(89)) xor (A(51) and B(88)) xor (A(52) and B(87)) xor (A(53) and B(86)) xor (A(54) and B(85)) xor (A(55) and B(84)) xor (A(56) and B(83)) xor (A(57) and B(82)) xor (A(58) and B(81)) xor (A(59) and B(80)) xor (A(60) and B(79)) xor (A(61) and B(78)) xor (A(62) and B(77)) xor (A(63) and B(76)) xor (A(64) and B(75)) xor (A(65) and B(74)) xor (A(66) and B(73)) xor (A(67) and B(72)) xor (A(68) and B(71)) xor (A(69) and B(70)) xor (A(70) and B(69)) xor (A(71) and B(68)) xor (A(72) and B(67)) xor (A(73) and B(66)) xor (A(74) and B(65)) xor (A(75) and B(64)) xor (A(76) and B(63)) xor (A(77) and B(62)) xor (A(78) and B(61)) xor (A(79) and B(60)) xor (A(80) and B(59)) xor (A(81) and B(58)) xor (A(82) and B(57)) xor (A(83) and B(56)) xor (A(84) and B(55)) xor (A(85) and B(54)) xor (A(86) and B(53)) xor (A(87) and B(52)) xor (A(88) and B(51)) xor (A(89) and B(50)) xor (A(90) and B(49)) xor (A(91) and B(48)) xor (A(92) and B(47)) xor (A(93) and B(46)) xor (A(94) and B(45)) xor (A(95) and B(44)) xor (A(96) and B(43)) xor (A(97) and B(42)) xor (A(98) and B(41)) xor (A(99) and B(40)) xor (A(100) and B(39)) xor (A(101) and B(38)) xor (A(102) and B(37)) xor (A(103) and B(36)) xor (A(104) and B(35)) xor (A(105) and B(34)) xor (A(106) and B(33)) xor (A(107) and B(32)) xor (A(108) and B(31)) xor (A(109) and B(30)) xor (A(110) and B(29)) xor (A(111) and B(28)) xor (A(112) and B(27)) xor (A(113) and B(26)) xor (A(114) and B(25)) xor (A(115) and B(24)) xor (A(116) and B(23)) xor (A(117) and B(23)) xor (A(118) and B(21)) xor (A(119) and B(20)) xor (A(120) and B(19)) xor (A(121) and B(18)) xor (A(122) and B(17)) xor (A(123) and B(16)) xor (A(124) and B(15)) xor (A(125) and B(14)) xor (A(126) and B(13)) xor (A(126) and B(127));
    C(13)  <= (A(0) and B(13)) xor (A(1) and B(12)) xor (A(2) and B(11)) xor (A(3) and B(10)) xor (A(4) and B(9)) xor (A(5) and B(8)) xor (A(6) and B(7)) xor (A(7) and B(6)) xor (A(8) and B(5)) xor (A(9) and B(4)) xor (A(10) and B(3)) xor (A(11) and B(2)) xor (A(12) and B(1)) xor (A(13) and B(0)) xor (A(6) and B(127)) xor (A(7) and B(126)) xor (A(8) and B(125)) xor (A(9) and B(124)) xor (A(10) and B(123)) xor (A(11) and B(122)) xor (A(12) and B(121)) xor (A(13) and B(120)) xor (A(14) and B(119)) xor (A(15) and B(118)) xor (A(16) and B(117)) xor (A(17) and B(116)) xor (A(18) and B(115)) xor (A(19) and B(114)) xor (A(20) and B(113)) xor (A(21) and B(112)) xor (A(23) and B(111)) xor (A(23) and B(110)) xor (A(24) and B(109)) xor (A(25) and B(108)) xor (A(26) and B(107)) xor (A(27) and B(106)) xor (A(28) and B(105)) xor (A(29) and B(104)) xor (A(30) and B(103)) xor (A(31) and B(102)) xor (A(32) and B(101)) xor (A(33) and B(100)) xor (A(34) and B(99)) xor (A(35) and B(98)) xor (A(36) and B(97)) xor (A(37) and B(96)) xor (A(38) and B(95)) xor (A(39) and B(94)) xor (A(40) and B(93)) xor (A(41) and B(92)) xor (A(42) and B(91)) xor (A(43) and B(90)) xor (A(44) and B(89)) xor (A(45) and B(88)) xor (A(46) and B(87)) xor (A(47) and B(86)) xor (A(48) and B(85)) xor (A(49) and B(84)) xor (A(50) and B(83)) xor (A(51) and B(82)) xor (A(52) and B(81)) xor (A(53) and B(80)) xor (A(54) and B(79)) xor (A(55) and B(78)) xor (A(56) and B(77)) xor (A(57) and B(76)) xor (A(58) and B(75)) xor (A(59) and B(74)) xor (A(60) and B(73)) xor (A(61) and B(72)) xor (A(62) and B(71)) xor (A(63) and B(70)) xor (A(64) and B(69)) xor (A(65) and B(68)) xor (A(66) and B(67)) xor (A(67) and B(66)) xor (A(68) and B(65)) xor (A(69) and B(64)) xor (A(70) and B(63)) xor (A(71) and B(62)) xor (A(72) and B(61)) xor (A(73) and B(60)) xor (A(74) and B(59)) xor (A(75) and B(58)) xor (A(76) and B(57)) xor (A(77) and B(56)) xor (A(78) and B(55)) xor (A(79) and B(54)) xor (A(80) and B(53)) xor (A(81) and B(52)) xor (A(82) and B(51)) xor (A(83) and B(50)) xor (A(84) and B(49)) xor (A(85) and B(48)) xor (A(86) and B(47)) xor (A(87) and B(46)) xor (A(88) and B(45)) xor (A(89) and B(44)) xor (A(90) and B(43)) xor (A(91) and B(42)) xor (A(92) and B(41)) xor (A(93) and B(40)) xor (A(94) and B(39)) xor (A(95) and B(38)) xor (A(96) and B(37)) xor (A(97) and B(36)) xor (A(98) and B(35)) xor (A(99) and B(34)) xor (A(100) and B(33)) xor (A(101) and B(32)) xor (A(102) and B(31)) xor (A(103) and B(30)) xor (A(104) and B(29)) xor (A(105) and B(28)) xor (A(106) and B(27)) xor (A(107) and B(26)) xor (A(108) and B(25)) xor (A(109) and B(24)) xor (A(110) and B(23)) xor (A(111) and B(23)) xor (A(112) and B(21)) xor (A(113) and B(20)) xor (A(114) and B(19)) xor (A(115) and B(18)) xor (A(116) and B(17)) xor (A(117) and B(16)) xor (A(118) and B(15)) xor (A(119) and B(14)) xor (A(120) and B(13)) xor (A(121) and B(12)) xor (A(122) and B(11)) xor (A(123) and B(10)) xor (A(124) and B(9)) xor (A(125) and B(8)) xor (A(126) and B(7)) xor (A(11) and B(127)) xor (A(12) and B(126)) xor (A(13) and B(125)) xor (A(14) and B(124)) xor (A(15) and B(123)) xor (A(16) and B(122)) xor (A(17) and B(121)) xor (A(18) and B(120)) xor (A(19) and B(119)) xor (A(20) and B(118)) xor (A(21) and B(117)) xor (A(23) and B(116)) xor (A(23) and B(115)) xor (A(24) and B(114)) xor (A(25) and B(113)) xor (A(26) and B(112)) xor (A(27) and B(111)) xor (A(28) and B(110)) xor (A(29) and B(109)) xor (A(30) and B(108)) xor (A(31) and B(107)) xor (A(32) and B(106)) xor (A(33) and B(105)) xor (A(34) and B(104)) xor (A(35) and B(103)) xor (A(36) and B(102)) xor (A(37) and B(101)) xor (A(38) and B(100)) xor (A(39) and B(99)) xor (A(40) and B(98)) xor (A(41) and B(97)) xor (A(42) and B(96)) xor (A(43) and B(95)) xor (A(44) and B(94)) xor (A(45) and B(93)) xor (A(46) and B(92)) xor (A(47) and B(91)) xor (A(48) and B(90)) xor (A(49) and B(89)) xor (A(50) and B(88)) xor (A(51) and B(87)) xor (A(52) and B(86)) xor (A(53) and B(85)) xor (A(54) and B(84)) xor (A(55) and B(83)) xor (A(56) and B(82)) xor (A(57) and B(81)) xor (A(58) and B(80)) xor (A(59) and B(79)) xor (A(60) and B(78)) xor (A(61) and B(77)) xor (A(62) and B(76)) xor (A(63) and B(75)) xor (A(64) and B(74)) xor (A(65) and B(73)) xor (A(66) and B(72)) xor (A(67) and B(71)) xor (A(68) and B(70)) xor (A(69) and B(69)) xor (A(70) and B(68)) xor (A(71) and B(67)) xor (A(72) and B(66)) xor (A(73) and B(65)) xor (A(74) and B(64)) xor (A(75) and B(63)) xor (A(76) and B(62)) xor (A(77) and B(61)) xor (A(78) and B(60)) xor (A(79) and B(59)) xor (A(80) and B(58)) xor (A(81) and B(57)) xor (A(82) and B(56)) xor (A(83) and B(55)) xor (A(84) and B(54)) xor (A(85) and B(53)) xor (A(86) and B(52)) xor (A(87) and B(51)) xor (A(88) and B(50)) xor (A(89) and B(49)) xor (A(90) and B(48)) xor (A(91) and B(47)) xor (A(92) and B(46)) xor (A(93) and B(45)) xor (A(94) and B(44)) xor (A(95) and B(43)) xor (A(96) and B(42)) xor (A(97) and B(41)) xor (A(98) and B(40)) xor (A(99) and B(39)) xor (A(100) and B(38)) xor (A(101) and B(37)) xor (A(102) and B(36)) xor (A(103) and B(35)) xor (A(104) and B(34)) xor (A(105) and B(33)) xor (A(106) and B(32)) xor (A(107) and B(31)) xor (A(108) and B(30)) xor (A(109) and B(29)) xor (A(110) and B(28)) xor (A(111) and B(27)) xor (A(112) and B(26)) xor (A(113) and B(25)) xor (A(114) and B(24)) xor (A(115) and B(23)) xor (A(116) and B(23)) xor (A(117) and B(21)) xor (A(118) and B(20)) xor (A(119) and B(19)) xor (A(120) and B(18)) xor (A(121) and B(17)) xor (A(122) and B(16)) xor (A(123) and B(15)) xor (A(124) and B(14)) xor (A(125) and B(13)) xor (A(126) and B(12)) xor (A(12) and B(127)) xor (A(13) and B(126)) xor (A(14) and B(125)) xor (A(15) and B(124)) xor (A(16) and B(123)) xor (A(17) and B(122)) xor (A(18) and B(121)) xor (A(19) and B(120)) xor (A(20) and B(119)) xor (A(21) and B(118)) xor (A(23) and B(117)) xor (A(23) and B(116)) xor (A(24) and B(115)) xor (A(25) and B(114)) xor (A(26) and B(113)) xor (A(27) and B(112)) xor (A(28) and B(111)) xor (A(29) and B(110)) xor (A(30) and B(109)) xor (A(31) and B(108)) xor (A(32) and B(107)) xor (A(33) and B(106)) xor (A(34) and B(105)) xor (A(35) and B(104)) xor (A(36) and B(103)) xor (A(37) and B(102)) xor (A(38) and B(101)) xor (A(39) and B(100)) xor (A(40) and B(99)) xor (A(41) and B(98)) xor (A(42) and B(97)) xor (A(43) and B(96)) xor (A(44) and B(95)) xor (A(45) and B(94)) xor (A(46) and B(93)) xor (A(47) and B(92)) xor (A(48) and B(91)) xor (A(49) and B(90)) xor (A(50) and B(89)) xor (A(51) and B(88)) xor (A(52) and B(87)) xor (A(53) and B(86)) xor (A(54) and B(85)) xor (A(55) and B(84)) xor (A(56) and B(83)) xor (A(57) and B(82)) xor (A(58) and B(81)) xor (A(59) and B(80)) xor (A(60) and B(79)) xor (A(61) and B(78)) xor (A(62) and B(77)) xor (A(63) and B(76)) xor (A(64) and B(75)) xor (A(65) and B(74)) xor (A(66) and B(73)) xor (A(67) and B(72)) xor (A(68) and B(71)) xor (A(69) and B(70)) xor (A(70) and B(69)) xor (A(71) and B(68)) xor (A(72) and B(67)) xor (A(73) and B(66)) xor (A(74) and B(65)) xor (A(75) and B(64)) xor (A(76) and B(63)) xor (A(77) and B(62)) xor (A(78) and B(61)) xor (A(79) and B(60)) xor (A(80) and B(59)) xor (A(81) and B(58)) xor (A(82) and B(57)) xor (A(83) and B(56)) xor (A(84) and B(55)) xor (A(85) and B(54)) xor (A(86) and B(53)) xor (A(87) and B(52)) xor (A(88) and B(51)) xor (A(89) and B(50)) xor (A(90) and B(49)) xor (A(91) and B(48)) xor (A(92) and B(47)) xor (A(93) and B(46)) xor (A(94) and B(45)) xor (A(95) and B(44)) xor (A(96) and B(43)) xor (A(97) and B(42)) xor (A(98) and B(41)) xor (A(99) and B(40)) xor (A(100) and B(39)) xor (A(101) and B(38)) xor (A(102) and B(37)) xor (A(103) and B(36)) xor (A(104) and B(35)) xor (A(105) and B(34)) xor (A(106) and B(33)) xor (A(107) and B(32)) xor (A(108) and B(31)) xor (A(109) and B(30)) xor (A(110) and B(29)) xor (A(111) and B(28)) xor (A(112) and B(27)) xor (A(113) and B(26)) xor (A(114) and B(25)) xor (A(115) and B(24)) xor (A(116) and B(23)) xor (A(117) and B(23)) xor (A(118) and B(21)) xor (A(119) and B(20)) xor (A(120) and B(19)) xor (A(121) and B(18)) xor (A(122) and B(17)) xor (A(123) and B(16)) xor (A(124) and B(15)) xor (A(125) and B(14)) xor (A(126) and B(13)) xor (A(13) and B(127)) xor (A(14) and B(126)) xor (A(15) and B(125)) xor (A(16) and B(124)) xor (A(17) and B(123)) xor (A(18) and B(122)) xor (A(19) and B(121)) xor (A(20) and B(120)) xor (A(21) and B(119)) xor (A(23) and B(118)) xor (A(23) and B(117)) xor (A(24) and B(116)) xor (A(25) and B(115)) xor (A(26) and B(114)) xor (A(27) and B(113)) xor (A(28) and B(112)) xor (A(29) and B(111)) xor (A(30) and B(110)) xor (A(31) and B(109)) xor (A(32) and B(108)) xor (A(33) and B(107)) xor (A(34) and B(106)) xor (A(35) and B(105)) xor (A(36) and B(104)) xor (A(37) and B(103)) xor (A(38) and B(102)) xor (A(39) and B(101)) xor (A(40) and B(100)) xor (A(41) and B(99)) xor (A(42) and B(98)) xor (A(43) and B(97)) xor (A(44) and B(96)) xor (A(45) and B(95)) xor (A(46) and B(94)) xor (A(47) and B(93)) xor (A(48) and B(92)) xor (A(49) and B(91)) xor (A(50) and B(90)) xor (A(51) and B(89)) xor (A(52) and B(88)) xor (A(53) and B(87)) xor (A(54) and B(86)) xor (A(55) and B(85)) xor (A(56) and B(84)) xor (A(57) and B(83)) xor (A(58) and B(82)) xor (A(59) and B(81)) xor (A(60) and B(80)) xor (A(61) and B(79)) xor (A(62) and B(78)) xor (A(63) and B(77)) xor (A(64) and B(76)) xor (A(65) and B(75)) xor (A(66) and B(74)) xor (A(67) and B(73)) xor (A(68) and B(72)) xor (A(69) and B(71)) xor (A(70) and B(70)) xor (A(71) and B(69)) xor (A(72) and B(68)) xor (A(73) and B(67)) xor (A(74) and B(66)) xor (A(75) and B(65)) xor (A(76) and B(64)) xor (A(77) and B(63)) xor (A(78) and B(62)) xor (A(79) and B(61)) xor (A(80) and B(60)) xor (A(81) and B(59)) xor (A(82) and B(58)) xor (A(83) and B(57)) xor (A(84) and B(56)) xor (A(85) and B(55)) xor (A(86) and B(54)) xor (A(87) and B(53)) xor (A(88) and B(52)) xor (A(89) and B(51)) xor (A(90) and B(50)) xor (A(91) and B(49)) xor (A(92) and B(48)) xor (A(93) and B(47)) xor (A(94) and B(46)) xor (A(95) and B(45)) xor (A(96) and B(44)) xor (A(97) and B(43)) xor (A(98) and B(42)) xor (A(99) and B(41)) xor (A(100) and B(40)) xor (A(101) and B(39)) xor (A(102) and B(38)) xor (A(103) and B(37)) xor (A(104) and B(36)) xor (A(105) and B(35)) xor (A(106) and B(34)) xor (A(107) and B(33)) xor (A(108) and B(32)) xor (A(109) and B(31)) xor (A(110) and B(30)) xor (A(111) and B(29)) xor (A(112) and B(28)) xor (A(113) and B(27)) xor (A(114) and B(26)) xor (A(115) and B(25)) xor (A(116) and B(24)) xor (A(117) and B(23)) xor (A(118) and B(23)) xor (A(119) and B(21)) xor (A(120) and B(20)) xor (A(121) and B(19)) xor (A(122) and B(18)) xor (A(123) and B(17)) xor (A(124) and B(16)) xor (A(125) and B(15)) xor (A(126) and B(15));
    C(14)  <= (A(0) and B(14)) xor (A(1) and B(13)) xor (A(2) and B(12)) xor (A(3) and B(11)) xor (A(4) and B(10)) xor (A(5) and B(9)) xor (A(6) and B(8)) xor (A(7) and B(7)) xor (A(8) and B(6)) xor (A(9) and B(5)) xor (A(10) and B(4)) xor (A(11) and B(3)) xor (A(12) and B(2)) xor (A(13) and B(1)) xor (A(14) and B(0)) xor (A(7) and B(127)) xor (A(8) and B(126)) xor (A(9) and B(125)) xor (A(10) and B(124)) xor (A(11) and B(123)) xor (A(12) and B(122)) xor (A(13) and B(121)) xor (A(14) and B(120)) xor (A(15) and B(119)) xor (A(16) and B(118)) xor (A(17) and B(117)) xor (A(18) and B(116)) xor (A(19) and B(115)) xor (A(20) and B(114)) xor (A(21) and B(113)) xor (A(23) and B(112)) xor (A(23) and B(111)) xor (A(24) and B(110)) xor (A(25) and B(109)) xor (A(26) and B(108)) xor (A(27) and B(107)) xor (A(28) and B(106)) xor (A(29) and B(105)) xor (A(30) and B(104)) xor (A(31) and B(103)) xor (A(32) and B(102)) xor (A(33) and B(101)) xor (A(34) and B(100)) xor (A(35) and B(99)) xor (A(36) and B(98)) xor (A(37) and B(97)) xor (A(38) and B(96)) xor (A(39) and B(95)) xor (A(40) and B(94)) xor (A(41) and B(93)) xor (A(42) and B(92)) xor (A(43) and B(91)) xor (A(44) and B(90)) xor (A(45) and B(89)) xor (A(46) and B(88)) xor (A(47) and B(87)) xor (A(48) and B(86)) xor (A(49) and B(85)) xor (A(50) and B(84)) xor (A(51) and B(83)) xor (A(52) and B(82)) xor (A(53) and B(81)) xor (A(54) and B(80)) xor (A(55) and B(79)) xor (A(56) and B(78)) xor (A(57) and B(77)) xor (A(58) and B(76)) xor (A(59) and B(75)) xor (A(60) and B(74)) xor (A(61) and B(73)) xor (A(62) and B(72)) xor (A(63) and B(71)) xor (A(64) and B(70)) xor (A(65) and B(69)) xor (A(66) and B(68)) xor (A(67) and B(67)) xor (A(68) and B(66)) xor (A(69) and B(65)) xor (A(70) and B(64)) xor (A(71) and B(63)) xor (A(72) and B(62)) xor (A(73) and B(61)) xor (A(74) and B(60)) xor (A(75) and B(59)) xor (A(76) and B(58)) xor (A(77) and B(57)) xor (A(78) and B(56)) xor (A(79) and B(55)) xor (A(80) and B(54)) xor (A(81) and B(53)) xor (A(82) and B(52)) xor (A(83) and B(51)) xor (A(84) and B(50)) xor (A(85) and B(49)) xor (A(86) and B(48)) xor (A(87) and B(47)) xor (A(88) and B(46)) xor (A(89) and B(45)) xor (A(90) and B(44)) xor (A(91) and B(43)) xor (A(92) and B(42)) xor (A(93) and B(41)) xor (A(94) and B(40)) xor (A(95) and B(39)) xor (A(96) and B(38)) xor (A(97) and B(37)) xor (A(98) and B(36)) xor (A(99) and B(35)) xor (A(100) and B(34)) xor (A(101) and B(33)) xor (A(102) and B(32)) xor (A(103) and B(31)) xor (A(104) and B(30)) xor (A(105) and B(29)) xor (A(106) and B(28)) xor (A(107) and B(27)) xor (A(108) and B(26)) xor (A(109) and B(25)) xor (A(110) and B(24)) xor (A(111) and B(23)) xor (A(112) and B(23)) xor (A(113) and B(21)) xor (A(114) and B(20)) xor (A(115) and B(19)) xor (A(116) and B(18)) xor (A(117) and B(17)) xor (A(118) and B(16)) xor (A(119) and B(15)) xor (A(120) and B(14)) xor (A(121) and B(13)) xor (A(122) and B(12)) xor (A(123) and B(11)) xor (A(124) and B(10)) xor (A(125) and B(9)) xor (A(126) and B(8)) xor (A(12) and B(127)) xor (A(13) and B(126)) xor (A(14) and B(125)) xor (A(15) and B(124)) xor (A(16) and B(123)) xor (A(17) and B(122)) xor (A(18) and B(121)) xor (A(19) and B(120)) xor (A(20) and B(119)) xor (A(21) and B(118)) xor (A(23) and B(117)) xor (A(23) and B(116)) xor (A(24) and B(115)) xor (A(25) and B(114)) xor (A(26) and B(113)) xor (A(27) and B(112)) xor (A(28) and B(111)) xor (A(29) and B(110)) xor (A(30) and B(109)) xor (A(31) and B(108)) xor (A(32) and B(107)) xor (A(33) and B(106)) xor (A(34) and B(105)) xor (A(35) and B(104)) xor (A(36) and B(103)) xor (A(37) and B(102)) xor (A(38) and B(101)) xor (A(39) and B(100)) xor (A(40) and B(99)) xor (A(41) and B(98)) xor (A(42) and B(97)) xor (A(43) and B(96)) xor (A(44) and B(95)) xor (A(45) and B(94)) xor (A(46) and B(93)) xor (A(47) and B(92)) xor (A(48) and B(91)) xor (A(49) and B(90)) xor (A(50) and B(89)) xor (A(51) and B(88)) xor (A(52) and B(87)) xor (A(53) and B(86)) xor (A(54) and B(85)) xor (A(55) and B(84)) xor (A(56) and B(83)) xor (A(57) and B(82)) xor (A(58) and B(81)) xor (A(59) and B(80)) xor (A(60) and B(79)) xor (A(61) and B(78)) xor (A(62) and B(77)) xor (A(63) and B(76)) xor (A(64) and B(75)) xor (A(65) and B(74)) xor (A(66) and B(73)) xor (A(67) and B(72)) xor (A(68) and B(71)) xor (A(69) and B(70)) xor (A(70) and B(69)) xor (A(71) and B(68)) xor (A(72) and B(67)) xor (A(73) and B(66)) xor (A(74) and B(65)) xor (A(75) and B(64)) xor (A(76) and B(63)) xor (A(77) and B(62)) xor (A(78) and B(61)) xor (A(79) and B(60)) xor (A(80) and B(59)) xor (A(81) and B(58)) xor (A(82) and B(57)) xor (A(83) and B(56)) xor (A(84) and B(55)) xor (A(85) and B(54)) xor (A(86) and B(53)) xor (A(87) and B(52)) xor (A(88) and B(51)) xor (A(89) and B(50)) xor (A(90) and B(49)) xor (A(91) and B(48)) xor (A(92) and B(47)) xor (A(93) and B(46)) xor (A(94) and B(45)) xor (A(95) and B(44)) xor (A(96) and B(43)) xor (A(97) and B(42)) xor (A(98) and B(41)) xor (A(99) and B(40)) xor (A(100) and B(39)) xor (A(101) and B(38)) xor (A(102) and B(37)) xor (A(103) and B(36)) xor (A(104) and B(35)) xor (A(105) and B(34)) xor (A(106) and B(33)) xor (A(107) and B(32)) xor (A(108) and B(31)) xor (A(109) and B(30)) xor (A(110) and B(29)) xor (A(111) and B(28)) xor (A(112) and B(27)) xor (A(113) and B(26)) xor (A(114) and B(25)) xor (A(115) and B(24)) xor (A(116) and B(23)) xor (A(117) and B(23)) xor (A(118) and B(21)) xor (A(119) and B(20)) xor (A(120) and B(19)) xor (A(121) and B(18)) xor (A(122) and B(17)) xor (A(123) and B(16)) xor (A(124) and B(15)) xor (A(125) and B(14)) xor (A(126) and B(13)) xor (A(13) and B(127)) xor (A(14) and B(126)) xor (A(15) and B(125)) xor (A(16) and B(124)) xor (A(17) and B(123)) xor (A(18) and B(122)) xor (A(19) and B(121)) xor (A(20) and B(120)) xor (A(21) and B(119)) xor (A(23) and B(118)) xor (A(23) and B(117)) xor (A(24) and B(116)) xor (A(25) and B(115)) xor (A(26) and B(114)) xor (A(27) and B(113)) xor (A(28) and B(112)) xor (A(29) and B(111)) xor (A(30) and B(110)) xor (A(31) and B(109)) xor (A(32) and B(108)) xor (A(33) and B(107)) xor (A(34) and B(106)) xor (A(35) and B(105)) xor (A(36) and B(104)) xor (A(37) and B(103)) xor (A(38) and B(102)) xor (A(39) and B(101)) xor (A(40) and B(100)) xor (A(41) and B(99)) xor (A(42) and B(98)) xor (A(43) and B(97)) xor (A(44) and B(96)) xor (A(45) and B(95)) xor (A(46) and B(94)) xor (A(47) and B(93)) xor (A(48) and B(92)) xor (A(49) and B(91)) xor (A(50) and B(90)) xor (A(51) and B(89)) xor (A(52) and B(88)) xor (A(53) and B(87)) xor (A(54) and B(86)) xor (A(55) and B(85)) xor (A(56) and B(84)) xor (A(57) and B(83)) xor (A(58) and B(82)) xor (A(59) and B(81)) xor (A(60) and B(80)) xor (A(61) and B(79)) xor (A(62) and B(78)) xor (A(63) and B(77)) xor (A(64) and B(76)) xor (A(65) and B(75)) xor (A(66) and B(74)) xor (A(67) and B(73)) xor (A(68) and B(72)) xor (A(69) and B(71)) xor (A(70) and B(70)) xor (A(71) and B(69)) xor (A(72) and B(68)) xor (A(73) and B(67)) xor (A(74) and B(66)) xor (A(75) and B(65)) xor (A(76) and B(64)) xor (A(77) and B(63)) xor (A(78) and B(62)) xor (A(79) and B(61)) xor (A(80) and B(60)) xor (A(81) and B(59)) xor (A(82) and B(58)) xor (A(83) and B(57)) xor (A(84) and B(56)) xor (A(85) and B(55)) xor (A(86) and B(54)) xor (A(87) and B(53)) xor (A(88) and B(52)) xor (A(89) and B(51)) xor (A(90) and B(50)) xor (A(91) and B(49)) xor (A(92) and B(48)) xor (A(93) and B(47)) xor (A(94) and B(46)) xor (A(95) and B(45)) xor (A(96) and B(44)) xor (A(97) and B(43)) xor (A(98) and B(42)) xor (A(99) and B(41)) xor (A(100) and B(40)) xor (A(101) and B(39)) xor (A(102) and B(38)) xor (A(103) and B(37)) xor (A(104) and B(36)) xor (A(105) and B(35)) xor (A(106) and B(34)) xor (A(107) and B(33)) xor (A(108) and B(32)) xor (A(109) and B(31)) xor (A(110) and B(30)) xor (A(111) and B(29)) xor (A(112) and B(28)) xor (A(113) and B(27)) xor (A(114) and B(26)) xor (A(115) and B(25)) xor (A(116) and B(24)) xor (A(117) and B(23)) xor (A(118) and B(23)) xor (A(119) and B(21)) xor (A(120) and B(20)) xor (A(121) and B(19)) xor (A(122) and B(18)) xor (A(123) and B(17)) xor (A(124) and B(16)) xor (A(125) and B(15)) xor (A(126) and B(14)) xor (A(14) and B(127)) xor (A(15) and B(126)) xor (A(16) and B(125)) xor (A(17) and B(124)) xor (A(18) and B(123)) xor (A(19) and B(122)) xor (A(20) and B(121)) xor (A(21) and B(120)) xor (A(23) and B(119)) xor (A(23) and B(118)) xor (A(24) and B(117)) xor (A(25) and B(116)) xor (A(26) and B(115)) xor (A(27) and B(114)) xor (A(28) and B(113)) xor (A(29) and B(112)) xor (A(30) and B(111)) xor (A(31) and B(110)) xor (A(32) and B(109)) xor (A(33) and B(108)) xor (A(34) and B(107)) xor (A(35) and B(106)) xor (A(36) and B(105)) xor (A(37) and B(104)) xor (A(38) and B(103)) xor (A(39) and B(102)) xor (A(40) and B(101)) xor (A(41) and B(100)) xor (A(42) and B(99)) xor (A(43) and B(98)) xor (A(44) and B(97)) xor (A(45) and B(96)) xor (A(46) and B(95)) xor (A(47) and B(94)) xor (A(48) and B(93)) xor (A(49) and B(92)) xor (A(50) and B(91)) xor (A(51) and B(90)) xor (A(52) and B(89)) xor (A(53) and B(88)) xor (A(54) and B(87)) xor (A(55) and B(86)) xor (A(56) and B(85)) xor (A(57) and B(84)) xor (A(58) and B(83)) xor (A(59) and B(82)) xor (A(60) and B(81)) xor (A(61) and B(80)) xor (A(62) and B(79)) xor (A(63) and B(78)) xor (A(64) and B(77)) xor (A(65) and B(76)) xor (A(66) and B(75)) xor (A(67) and B(74)) xor (A(68) and B(73)) xor (A(69) and B(72)) xor (A(70) and B(71)) xor (A(71) and B(70)) xor (A(72) and B(69)) xor (A(73) and B(68)) xor (A(74) and B(67)) xor (A(75) and B(66)) xor (A(76) and B(65)) xor (A(77) and B(64)) xor (A(78) and B(63)) xor (A(79) and B(62)) xor (A(80) and B(61)) xor (A(81) and B(60)) xor (A(82) and B(59)) xor (A(83) and B(58)) xor (A(84) and B(57)) xor (A(85) and B(56)) xor (A(86) and B(55)) xor (A(87) and B(54)) xor (A(88) and B(53)) xor (A(89) and B(52)) xor (A(90) and B(51)) xor (A(91) and B(50)) xor (A(92) and B(49)) xor (A(93) and B(48)) xor (A(94) and B(47)) xor (A(95) and B(46)) xor (A(96) and B(45)) xor (A(97) and B(44)) xor (A(98) and B(43)) xor (A(99) and B(42)) xor (A(100) and B(41)) xor (A(101) and B(40)) xor (A(102) and B(39)) xor (A(103) and B(38)) xor (A(104) and B(37)) xor (A(105) and B(36)) xor (A(106) and B(35)) xor (A(107) and B(34)) xor (A(108) and B(33)) xor (A(109) and B(32)) xor (A(110) and B(31)) xor (A(111) and B(30)) xor (A(112) and B(29)) xor (A(113) and B(28)) xor (A(114) and B(27)) xor (A(115) and B(26)) xor (A(116) and B(25)) xor (A(117) and B(24)) xor (A(118) and B(23)) xor (A(119) and B(23)) xor (A(120) and B(21)) xor (A(121) and B(20)) xor (A(122) and B(19)) xor (A(123) and B(18)) xor (A(124) and B(17)) xor (A(125) and B(16)) xor (A(126) and B(16));
    C(15)  <= (A(0) and B(15)) xor (A(1) and B(14)) xor (A(2) and B(13)) xor (A(3) and B(12)) xor (A(4) and B(11)) xor (A(5) and B(10)) xor (A(6) and B(9)) xor (A(7) and B(8)) xor (A(8) and B(7)) xor (A(9) and B(6)) xor (A(10) and B(5)) xor (A(11) and B(4)) xor (A(12) and B(3)) xor (A(13) and B(2)) xor (A(14) and B(1)) xor (A(15) and B(0)) xor (A(8) and B(127)) xor (A(9) and B(126)) xor (A(10) and B(125)) xor (A(11) and B(124)) xor (A(12) and B(123)) xor (A(13) and B(122)) xor (A(14) and B(121)) xor (A(15) and B(120)) xor (A(16) and B(119)) xor (A(17) and B(118)) xor (A(18) and B(117)) xor (A(19) and B(116)) xor (A(20) and B(115)) xor (A(21) and B(114)) xor (A(23) and B(113)) xor (A(23) and B(112)) xor (A(24) and B(111)) xor (A(25) and B(110)) xor (A(26) and B(109)) xor (A(27) and B(108)) xor (A(28) and B(107)) xor (A(29) and B(106)) xor (A(30) and B(105)) xor (A(31) and B(104)) xor (A(32) and B(103)) xor (A(33) and B(102)) xor (A(34) and B(101)) xor (A(35) and B(100)) xor (A(36) and B(99)) xor (A(37) and B(98)) xor (A(38) and B(97)) xor (A(39) and B(96)) xor (A(40) and B(95)) xor (A(41) and B(94)) xor (A(42) and B(93)) xor (A(43) and B(92)) xor (A(44) and B(91)) xor (A(45) and B(90)) xor (A(46) and B(89)) xor (A(47) and B(88)) xor (A(48) and B(87)) xor (A(49) and B(86)) xor (A(50) and B(85)) xor (A(51) and B(84)) xor (A(52) and B(83)) xor (A(53) and B(82)) xor (A(54) and B(81)) xor (A(55) and B(80)) xor (A(56) and B(79)) xor (A(57) and B(78)) xor (A(58) and B(77)) xor (A(59) and B(76)) xor (A(60) and B(75)) xor (A(61) and B(74)) xor (A(62) and B(73)) xor (A(63) and B(72)) xor (A(64) and B(71)) xor (A(65) and B(70)) xor (A(66) and B(69)) xor (A(67) and B(68)) xor (A(68) and B(67)) xor (A(69) and B(66)) xor (A(70) and B(65)) xor (A(71) and B(64)) xor (A(72) and B(63)) xor (A(73) and B(62)) xor (A(74) and B(61)) xor (A(75) and B(60)) xor (A(76) and B(59)) xor (A(77) and B(58)) xor (A(78) and B(57)) xor (A(79) and B(56)) xor (A(80) and B(55)) xor (A(81) and B(54)) xor (A(82) and B(53)) xor (A(83) and B(52)) xor (A(84) and B(51)) xor (A(85) and B(50)) xor (A(86) and B(49)) xor (A(87) and B(48)) xor (A(88) and B(47)) xor (A(89) and B(46)) xor (A(90) and B(45)) xor (A(91) and B(44)) xor (A(92) and B(43)) xor (A(93) and B(42)) xor (A(94) and B(41)) xor (A(95) and B(40)) xor (A(96) and B(39)) xor (A(97) and B(38)) xor (A(98) and B(37)) xor (A(99) and B(36)) xor (A(100) and B(35)) xor (A(101) and B(34)) xor (A(102) and B(33)) xor (A(103) and B(32)) xor (A(104) and B(31)) xor (A(105) and B(30)) xor (A(106) and B(29)) xor (A(107) and B(28)) xor (A(108) and B(27)) xor (A(109) and B(26)) xor (A(110) and B(25)) xor (A(111) and B(24)) xor (A(112) and B(23)) xor (A(113) and B(23)) xor (A(114) and B(21)) xor (A(115) and B(20)) xor (A(116) and B(19)) xor (A(117) and B(18)) xor (A(118) and B(17)) xor (A(119) and B(16)) xor (A(120) and B(15)) xor (A(121) and B(14)) xor (A(122) and B(13)) xor (A(123) and B(12)) xor (A(124) and B(11)) xor (A(125) and B(10)) xor (A(126) and B(9)) xor (A(13) and B(127)) xor (A(14) and B(126)) xor (A(15) and B(125)) xor (A(16) and B(124)) xor (A(17) and B(123)) xor (A(18) and B(122)) xor (A(19) and B(121)) xor (A(20) and B(120)) xor (A(21) and B(119)) xor (A(23) and B(118)) xor (A(23) and B(117)) xor (A(24) and B(116)) xor (A(25) and B(115)) xor (A(26) and B(114)) xor (A(27) and B(113)) xor (A(28) and B(112)) xor (A(29) and B(111)) xor (A(30) and B(110)) xor (A(31) and B(109)) xor (A(32) and B(108)) xor (A(33) and B(107)) xor (A(34) and B(106)) xor (A(35) and B(105)) xor (A(36) and B(104)) xor (A(37) and B(103)) xor (A(38) and B(102)) xor (A(39) and B(101)) xor (A(40) and B(100)) xor (A(41) and B(99)) xor (A(42) and B(98)) xor (A(43) and B(97)) xor (A(44) and B(96)) xor (A(45) and B(95)) xor (A(46) and B(94)) xor (A(47) and B(93)) xor (A(48) and B(92)) xor (A(49) and B(91)) xor (A(50) and B(90)) xor (A(51) and B(89)) xor (A(52) and B(88)) xor (A(53) and B(87)) xor (A(54) and B(86)) xor (A(55) and B(85)) xor (A(56) and B(84)) xor (A(57) and B(83)) xor (A(58) and B(82)) xor (A(59) and B(81)) xor (A(60) and B(80)) xor (A(61) and B(79)) xor (A(62) and B(78)) xor (A(63) and B(77)) xor (A(64) and B(76)) xor (A(65) and B(75)) xor (A(66) and B(74)) xor (A(67) and B(73)) xor (A(68) and B(72)) xor (A(69) and B(71)) xor (A(70) and B(70)) xor (A(71) and B(69)) xor (A(72) and B(68)) xor (A(73) and B(67)) xor (A(74) and B(66)) xor (A(75) and B(65)) xor (A(76) and B(64)) xor (A(77) and B(63)) xor (A(78) and B(62)) xor (A(79) and B(61)) xor (A(80) and B(60)) xor (A(81) and B(59)) xor (A(82) and B(58)) xor (A(83) and B(57)) xor (A(84) and B(56)) xor (A(85) and B(55)) xor (A(86) and B(54)) xor (A(87) and B(53)) xor (A(88) and B(52)) xor (A(89) and B(51)) xor (A(90) and B(50)) xor (A(91) and B(49)) xor (A(92) and B(48)) xor (A(93) and B(47)) xor (A(94) and B(46)) xor (A(95) and B(45)) xor (A(96) and B(44)) xor (A(97) and B(43)) xor (A(98) and B(42)) xor (A(99) and B(41)) xor (A(100) and B(40)) xor (A(101) and B(39)) xor (A(102) and B(38)) xor (A(103) and B(37)) xor (A(104) and B(36)) xor (A(105) and B(35)) xor (A(106) and B(34)) xor (A(107) and B(33)) xor (A(108) and B(32)) xor (A(109) and B(31)) xor (A(110) and B(30)) xor (A(111) and B(29)) xor (A(112) and B(28)) xor (A(113) and B(27)) xor (A(114) and B(26)) xor (A(115) and B(25)) xor (A(116) and B(24)) xor (A(117) and B(23)) xor (A(118) and B(23)) xor (A(119) and B(21)) xor (A(120) and B(20)) xor (A(121) and B(19)) xor (A(122) and B(18)) xor (A(123) and B(17)) xor (A(124) and B(16)) xor (A(125) and B(15)) xor (A(126) and B(14)) xor (A(14) and B(127)) xor (A(15) and B(126)) xor (A(16) and B(125)) xor (A(17) and B(124)) xor (A(18) and B(123)) xor (A(19) and B(122)) xor (A(20) and B(121)) xor (A(21) and B(120)) xor (A(23) and B(119)) xor (A(23) and B(118)) xor (A(24) and B(117)) xor (A(25) and B(116)) xor (A(26) and B(115)) xor (A(27) and B(114)) xor (A(28) and B(113)) xor (A(29) and B(112)) xor (A(30) and B(111)) xor (A(31) and B(110)) xor (A(32) and B(109)) xor (A(33) and B(108)) xor (A(34) and B(107)) xor (A(35) and B(106)) xor (A(36) and B(105)) xor (A(37) and B(104)) xor (A(38) and B(103)) xor (A(39) and B(102)) xor (A(40) and B(101)) xor (A(41) and B(100)) xor (A(42) and B(99)) xor (A(43) and B(98)) xor (A(44) and B(97)) xor (A(45) and B(96)) xor (A(46) and B(95)) xor (A(47) and B(94)) xor (A(48) and B(93)) xor (A(49) and B(92)) xor (A(50) and B(91)) xor (A(51) and B(90)) xor (A(52) and B(89)) xor (A(53) and B(88)) xor (A(54) and B(87)) xor (A(55) and B(86)) xor (A(56) and B(85)) xor (A(57) and B(84)) xor (A(58) and B(83)) xor (A(59) and B(82)) xor (A(60) and B(81)) xor (A(61) and B(80)) xor (A(62) and B(79)) xor (A(63) and B(78)) xor (A(64) and B(77)) xor (A(65) and B(76)) xor (A(66) and B(75)) xor (A(67) and B(74)) xor (A(68) and B(73)) xor (A(69) and B(72)) xor (A(70) and B(71)) xor (A(71) and B(70)) xor (A(72) and B(69)) xor (A(73) and B(68)) xor (A(74) and B(67)) xor (A(75) and B(66)) xor (A(76) and B(65)) xor (A(77) and B(64)) xor (A(78) and B(63)) xor (A(79) and B(62)) xor (A(80) and B(61)) xor (A(81) and B(60)) xor (A(82) and B(59)) xor (A(83) and B(58)) xor (A(84) and B(57)) xor (A(85) and B(56)) xor (A(86) and B(55)) xor (A(87) and B(54)) xor (A(88) and B(53)) xor (A(89) and B(52)) xor (A(90) and B(51)) xor (A(91) and B(50)) xor (A(92) and B(49)) xor (A(93) and B(48)) xor (A(94) and B(47)) xor (A(95) and B(46)) xor (A(96) and B(45)) xor (A(97) and B(44)) xor (A(98) and B(43)) xor (A(99) and B(42)) xor (A(100) and B(41)) xor (A(101) and B(40)) xor (A(102) and B(39)) xor (A(103) and B(38)) xor (A(104) and B(37)) xor (A(105) and B(36)) xor (A(106) and B(35)) xor (A(107) and B(34)) xor (A(108) and B(33)) xor (A(109) and B(32)) xor (A(110) and B(31)) xor (A(111) and B(30)) xor (A(112) and B(29)) xor (A(113) and B(28)) xor (A(114) and B(27)) xor (A(115) and B(26)) xor (A(116) and B(25)) xor (A(117) and B(24)) xor (A(118) and B(23)) xor (A(119) and B(23)) xor (A(120) and B(21)) xor (A(121) and B(20)) xor (A(122) and B(19)) xor (A(123) and B(18)) xor (A(124) and B(17)) xor (A(125) and B(16)) xor (A(126) and B(15)) xor (A(15) and B(127)) xor (A(16) and B(126)) xor (A(17) and B(125)) xor (A(18) and B(124)) xor (A(19) and B(123)) xor (A(20) and B(122)) xor (A(21) and B(121)) xor (A(23) and B(120)) xor (A(23) and B(119)) xor (A(24) and B(118)) xor (A(25) and B(117)) xor (A(26) and B(116)) xor (A(27) and B(115)) xor (A(28) and B(114)) xor (A(29) and B(113)) xor (A(30) and B(112)) xor (A(31) and B(111)) xor (A(32) and B(110)) xor (A(33) and B(109)) xor (A(34) and B(108)) xor (A(35) and B(107)) xor (A(36) and B(106)) xor (A(37) and B(105)) xor (A(38) and B(104)) xor (A(39) and B(103)) xor (A(40) and B(102)) xor (A(41) and B(101)) xor (A(42) and B(100)) xor (A(43) and B(99)) xor (A(44) and B(98)) xor (A(45) and B(97)) xor (A(46) and B(96)) xor (A(47) and B(95)) xor (A(48) and B(94)) xor (A(49) and B(93)) xor (A(50) and B(92)) xor (A(51) and B(91)) xor (A(52) and B(90)) xor (A(53) and B(89)) xor (A(54) and B(88)) xor (A(55) and B(87)) xor (A(56) and B(86)) xor (A(57) and B(85)) xor (A(58) and B(84)) xor (A(59) and B(83)) xor (A(60) and B(82)) xor (A(61) and B(81)) xor (A(62) and B(80)) xor (A(63) and B(79)) xor (A(64) and B(78)) xor (A(65) and B(77)) xor (A(66) and B(76)) xor (A(67) and B(75)) xor (A(68) and B(74)) xor (A(69) and B(73)) xor (A(70) and B(72)) xor (A(71) and B(71)) xor (A(72) and B(70)) xor (A(73) and B(69)) xor (A(74) and B(68)) xor (A(75) and B(67)) xor (A(76) and B(66)) xor (A(77) and B(65)) xor (A(78) and B(64)) xor (A(79) and B(63)) xor (A(80) and B(62)) xor (A(81) and B(61)) xor (A(82) and B(60)) xor (A(83) and B(59)) xor (A(84) and B(58)) xor (A(85) and B(57)) xor (A(86) and B(56)) xor (A(87) and B(55)) xor (A(88) and B(54)) xor (A(89) and B(53)) xor (A(90) and B(52)) xor (A(91) and B(51)) xor (A(92) and B(50)) xor (A(93) and B(49)) xor (A(94) and B(48)) xor (A(95) and B(47)) xor (A(96) and B(46)) xor (A(97) and B(45)) xor (A(98) and B(44)) xor (A(99) and B(43)) xor (A(100) and B(42)) xor (A(101) and B(41)) xor (A(102) and B(40)) xor (A(103) and B(39)) xor (A(104) and B(38)) xor (A(105) and B(37)) xor (A(106) and B(36)) xor (A(107) and B(35)) xor (A(108) and B(34)) xor (A(109) and B(33)) xor (A(110) and B(32)) xor (A(111) and B(31)) xor (A(112) and B(30)) xor (A(113) and B(29)) xor (A(114) and B(28)) xor (A(115) and B(27)) xor (A(116) and B(26)) xor (A(117) and B(25)) xor (A(118) and B(24)) xor (A(119) and B(23)) xor (A(120) and B(23)) xor (A(121) and B(21)) xor (A(122) and B(20)) xor (A(123) and B(19)) xor (A(124) and B(18)) xor (A(125) and B(17)) xor (A(126) and B(17));
    C(16)  <= (A(0) and B(16)) xor (A(1) and B(15)) xor (A(2) and B(14)) xor (A(3) and B(13)) xor (A(4) and B(12)) xor (A(5) and B(11)) xor (A(6) and B(10)) xor (A(7) and B(9)) xor (A(8) and B(8)) xor (A(9) and B(7)) xor (A(10) and B(6)) xor (A(11) and B(5)) xor (A(12) and B(4)) xor (A(13) and B(3)) xor (A(14) and B(2)) xor (A(15) and B(1)) xor (A(16) and B(0)) xor (A(9) and B(127)) xor (A(10) and B(126)) xor (A(11) and B(125)) xor (A(12) and B(124)) xor (A(13) and B(123)) xor (A(14) and B(122)) xor (A(15) and B(121)) xor (A(16) and B(120)) xor (A(17) and B(119)) xor (A(18) and B(118)) xor (A(19) and B(117)) xor (A(20) and B(116)) xor (A(21) and B(115)) xor (A(23) and B(114)) xor (A(23) and B(113)) xor (A(24) and B(112)) xor (A(25) and B(111)) xor (A(26) and B(110)) xor (A(27) and B(109)) xor (A(28) and B(108)) xor (A(29) and B(107)) xor (A(30) and B(106)) xor (A(31) and B(105)) xor (A(32) and B(104)) xor (A(33) and B(103)) xor (A(34) and B(102)) xor (A(35) and B(101)) xor (A(36) and B(100)) xor (A(37) and B(99)) xor (A(38) and B(98)) xor (A(39) and B(97)) xor (A(40) and B(96)) xor (A(41) and B(95)) xor (A(42) and B(94)) xor (A(43) and B(93)) xor (A(44) and B(92)) xor (A(45) and B(91)) xor (A(46) and B(90)) xor (A(47) and B(89)) xor (A(48) and B(88)) xor (A(49) and B(87)) xor (A(50) and B(86)) xor (A(51) and B(85)) xor (A(52) and B(84)) xor (A(53) and B(83)) xor (A(54) and B(82)) xor (A(55) and B(81)) xor (A(56) and B(80)) xor (A(57) and B(79)) xor (A(58) and B(78)) xor (A(59) and B(77)) xor (A(60) and B(76)) xor (A(61) and B(75)) xor (A(62) and B(74)) xor (A(63) and B(73)) xor (A(64) and B(72)) xor (A(65) and B(71)) xor (A(66) and B(70)) xor (A(67) and B(69)) xor (A(68) and B(68)) xor (A(69) and B(67)) xor (A(70) and B(66)) xor (A(71) and B(65)) xor (A(72) and B(64)) xor (A(73) and B(63)) xor (A(74) and B(62)) xor (A(75) and B(61)) xor (A(76) and B(60)) xor (A(77) and B(59)) xor (A(78) and B(58)) xor (A(79) and B(57)) xor (A(80) and B(56)) xor (A(81) and B(55)) xor (A(82) and B(54)) xor (A(83) and B(53)) xor (A(84) and B(52)) xor (A(85) and B(51)) xor (A(86) and B(50)) xor (A(87) and B(49)) xor (A(88) and B(48)) xor (A(89) and B(47)) xor (A(90) and B(46)) xor (A(91) and B(45)) xor (A(92) and B(44)) xor (A(93) and B(43)) xor (A(94) and B(42)) xor (A(95) and B(41)) xor (A(96) and B(40)) xor (A(97) and B(39)) xor (A(98) and B(38)) xor (A(99) and B(37)) xor (A(100) and B(36)) xor (A(101) and B(35)) xor (A(102) and B(34)) xor (A(103) and B(33)) xor (A(104) and B(32)) xor (A(105) and B(31)) xor (A(106) and B(30)) xor (A(107) and B(29)) xor (A(108) and B(28)) xor (A(109) and B(27)) xor (A(110) and B(26)) xor (A(111) and B(25)) xor (A(112) and B(24)) xor (A(113) and B(23)) xor (A(114) and B(23)) xor (A(115) and B(21)) xor (A(116) and B(20)) xor (A(117) and B(19)) xor (A(118) and B(18)) xor (A(119) and B(17)) xor (A(120) and B(16)) xor (A(121) and B(15)) xor (A(122) and B(14)) xor (A(123) and B(13)) xor (A(124) and B(12)) xor (A(125) and B(11)) xor (A(126) and B(10)) xor (A(14) and B(127)) xor (A(15) and B(126)) xor (A(16) and B(125)) xor (A(17) and B(124)) xor (A(18) and B(123)) xor (A(19) and B(122)) xor (A(20) and B(121)) xor (A(21) and B(120)) xor (A(23) and B(119)) xor (A(23) and B(118)) xor (A(24) and B(117)) xor (A(25) and B(116)) xor (A(26) and B(115)) xor (A(27) and B(114)) xor (A(28) and B(113)) xor (A(29) and B(112)) xor (A(30) and B(111)) xor (A(31) and B(110)) xor (A(32) and B(109)) xor (A(33) and B(108)) xor (A(34) and B(107)) xor (A(35) and B(106)) xor (A(36) and B(105)) xor (A(37) and B(104)) xor (A(38) and B(103)) xor (A(39) and B(102)) xor (A(40) and B(101)) xor (A(41) and B(100)) xor (A(42) and B(99)) xor (A(43) and B(98)) xor (A(44) and B(97)) xor (A(45) and B(96)) xor (A(46) and B(95)) xor (A(47) and B(94)) xor (A(48) and B(93)) xor (A(49) and B(92)) xor (A(50) and B(91)) xor (A(51) and B(90)) xor (A(52) and B(89)) xor (A(53) and B(88)) xor (A(54) and B(87)) xor (A(55) and B(86)) xor (A(56) and B(85)) xor (A(57) and B(84)) xor (A(58) and B(83)) xor (A(59) and B(82)) xor (A(60) and B(81)) xor (A(61) and B(80)) xor (A(62) and B(79)) xor (A(63) and B(78)) xor (A(64) and B(77)) xor (A(65) and B(76)) xor (A(66) and B(75)) xor (A(67) and B(74)) xor (A(68) and B(73)) xor (A(69) and B(72)) xor (A(70) and B(71)) xor (A(71) and B(70)) xor (A(72) and B(69)) xor (A(73) and B(68)) xor (A(74) and B(67)) xor (A(75) and B(66)) xor (A(76) and B(65)) xor (A(77) and B(64)) xor (A(78) and B(63)) xor (A(79) and B(62)) xor (A(80) and B(61)) xor (A(81) and B(60)) xor (A(82) and B(59)) xor (A(83) and B(58)) xor (A(84) and B(57)) xor (A(85) and B(56)) xor (A(86) and B(55)) xor (A(87) and B(54)) xor (A(88) and B(53)) xor (A(89) and B(52)) xor (A(90) and B(51)) xor (A(91) and B(50)) xor (A(92) and B(49)) xor (A(93) and B(48)) xor (A(94) and B(47)) xor (A(95) and B(46)) xor (A(96) and B(45)) xor (A(97) and B(44)) xor (A(98) and B(43)) xor (A(99) and B(42)) xor (A(100) and B(41)) xor (A(101) and B(40)) xor (A(102) and B(39)) xor (A(103) and B(38)) xor (A(104) and B(37)) xor (A(105) and B(36)) xor (A(106) and B(35)) xor (A(107) and B(34)) xor (A(108) and B(33)) xor (A(109) and B(32)) xor (A(110) and B(31)) xor (A(111) and B(30)) xor (A(112) and B(29)) xor (A(113) and B(28)) xor (A(114) and B(27)) xor (A(115) and B(26)) xor (A(116) and B(25)) xor (A(117) and B(24)) xor (A(118) and B(23)) xor (A(119) and B(23)) xor (A(120) and B(21)) xor (A(121) and B(20)) xor (A(122) and B(19)) xor (A(123) and B(18)) xor (A(124) and B(17)) xor (A(125) and B(16)) xor (A(126) and B(15)) xor (A(15) and B(127)) xor (A(16) and B(126)) xor (A(17) and B(125)) xor (A(18) and B(124)) xor (A(19) and B(123)) xor (A(20) and B(122)) xor (A(21) and B(121)) xor (A(23) and B(120)) xor (A(23) and B(119)) xor (A(24) and B(118)) xor (A(25) and B(117)) xor (A(26) and B(116)) xor (A(27) and B(115)) xor (A(28) and B(114)) xor (A(29) and B(113)) xor (A(30) and B(112)) xor (A(31) and B(111)) xor (A(32) and B(110)) xor (A(33) and B(109)) xor (A(34) and B(108)) xor (A(35) and B(107)) xor (A(36) and B(106)) xor (A(37) and B(105)) xor (A(38) and B(104)) xor (A(39) and B(103)) xor (A(40) and B(102)) xor (A(41) and B(101)) xor (A(42) and B(100)) xor (A(43) and B(99)) xor (A(44) and B(98)) xor (A(45) and B(97)) xor (A(46) and B(96)) xor (A(47) and B(95)) xor (A(48) and B(94)) xor (A(49) and B(93)) xor (A(50) and B(92)) xor (A(51) and B(91)) xor (A(52) and B(90)) xor (A(53) and B(89)) xor (A(54) and B(88)) xor (A(55) and B(87)) xor (A(56) and B(86)) xor (A(57) and B(85)) xor (A(58) and B(84)) xor (A(59) and B(83)) xor (A(60) and B(82)) xor (A(61) and B(81)) xor (A(62) and B(80)) xor (A(63) and B(79)) xor (A(64) and B(78)) xor (A(65) and B(77)) xor (A(66) and B(76)) xor (A(67) and B(75)) xor (A(68) and B(74)) xor (A(69) and B(73)) xor (A(70) and B(72)) xor (A(71) and B(71)) xor (A(72) and B(70)) xor (A(73) and B(69)) xor (A(74) and B(68)) xor (A(75) and B(67)) xor (A(76) and B(66)) xor (A(77) and B(65)) xor (A(78) and B(64)) xor (A(79) and B(63)) xor (A(80) and B(62)) xor (A(81) and B(61)) xor (A(82) and B(60)) xor (A(83) and B(59)) xor (A(84) and B(58)) xor (A(85) and B(57)) xor (A(86) and B(56)) xor (A(87) and B(55)) xor (A(88) and B(54)) xor (A(89) and B(53)) xor (A(90) and B(52)) xor (A(91) and B(51)) xor (A(92) and B(50)) xor (A(93) and B(49)) xor (A(94) and B(48)) xor (A(95) and B(47)) xor (A(96) and B(46)) xor (A(97) and B(45)) xor (A(98) and B(44)) xor (A(99) and B(43)) xor (A(100) and B(42)) xor (A(101) and B(41)) xor (A(102) and B(40)) xor (A(103) and B(39)) xor (A(104) and B(38)) xor (A(105) and B(37)) xor (A(106) and B(36)) xor (A(107) and B(35)) xor (A(108) and B(34)) xor (A(109) and B(33)) xor (A(110) and B(32)) xor (A(111) and B(31)) xor (A(112) and B(30)) xor (A(113) and B(29)) xor (A(114) and B(28)) xor (A(115) and B(27)) xor (A(116) and B(26)) xor (A(117) and B(25)) xor (A(118) and B(24)) xor (A(119) and B(23)) xor (A(120) and B(23)) xor (A(121) and B(21)) xor (A(122) and B(20)) xor (A(123) and B(19)) xor (A(124) and B(18)) xor (A(125) and B(17)) xor (A(126) and B(16)) xor (A(16) and B(127)) xor (A(17) and B(126)) xor (A(18) and B(125)) xor (A(19) and B(124)) xor (A(20) and B(123)) xor (A(21) and B(122)) xor (A(23) and B(121)) xor (A(23) and B(120)) xor (A(24) and B(119)) xor (A(25) and B(118)) xor (A(26) and B(117)) xor (A(27) and B(116)) xor (A(28) and B(115)) xor (A(29) and B(114)) xor (A(30) and B(113)) xor (A(31) and B(112)) xor (A(32) and B(111)) xor (A(33) and B(110)) xor (A(34) and B(109)) xor (A(35) and B(108)) xor (A(36) and B(107)) xor (A(37) and B(106)) xor (A(38) and B(105)) xor (A(39) and B(104)) xor (A(40) and B(103)) xor (A(41) and B(102)) xor (A(42) and B(101)) xor (A(43) and B(100)) xor (A(44) and B(99)) xor (A(45) and B(98)) xor (A(46) and B(97)) xor (A(47) and B(96)) xor (A(48) and B(95)) xor (A(49) and B(94)) xor (A(50) and B(93)) xor (A(51) and B(92)) xor (A(52) and B(91)) xor (A(53) and B(90)) xor (A(54) and B(89)) xor (A(55) and B(88)) xor (A(56) and B(87)) xor (A(57) and B(86)) xor (A(58) and B(85)) xor (A(59) and B(84)) xor (A(60) and B(83)) xor (A(61) and B(82)) xor (A(62) and B(81)) xor (A(63) and B(80)) xor (A(64) and B(79)) xor (A(65) and B(78)) xor (A(66) and B(77)) xor (A(67) and B(76)) xor (A(68) and B(75)) xor (A(69) and B(74)) xor (A(70) and B(73)) xor (A(71) and B(72)) xor (A(72) and B(71)) xor (A(73) and B(70)) xor (A(74) and B(69)) xor (A(75) and B(68)) xor (A(76) and B(67)) xor (A(77) and B(66)) xor (A(78) and B(65)) xor (A(79) and B(64)) xor (A(80) and B(63)) xor (A(81) and B(62)) xor (A(82) and B(61)) xor (A(83) and B(60)) xor (A(84) and B(59)) xor (A(85) and B(58)) xor (A(86) and B(57)) xor (A(87) and B(56)) xor (A(88) and B(55)) xor (A(89) and B(54)) xor (A(90) and B(53)) xor (A(91) and B(52)) xor (A(92) and B(51)) xor (A(93) and B(50)) xor (A(94) and B(49)) xor (A(95) and B(48)) xor (A(96) and B(47)) xor (A(97) and B(46)) xor (A(98) and B(45)) xor (A(99) and B(44)) xor (A(100) and B(43)) xor (A(101) and B(42)) xor (A(102) and B(41)) xor (A(103) and B(40)) xor (A(104) and B(39)) xor (A(105) and B(38)) xor (A(106) and B(37)) xor (A(107) and B(36)) xor (A(108) and B(35)) xor (A(109) and B(34)) xor (A(110) and B(33)) xor (A(111) and B(32)) xor (A(112) and B(31)) xor (A(113) and B(30)) xor (A(114) and B(29)) xor (A(115) and B(28)) xor (A(116) and B(27)) xor (A(117) and B(26)) xor (A(118) and B(25)) xor (A(119) and B(24)) xor (A(120) and B(23)) xor (A(121) and B(23)) xor (A(122) and B(21)) xor (A(123) and B(20)) xor (A(124) and B(19)) xor (A(125) and B(18)) xor (A(126) and B(18));
    C(17)  <= (A(0) and B(17)) xor (A(1) and B(16)) xor (A(2) and B(15)) xor (A(3) and B(14)) xor (A(4) and B(13)) xor (A(5) and B(12)) xor (A(6) and B(11)) xor (A(7) and B(10)) xor (A(8) and B(9)) xor (A(9) and B(8)) xor (A(10) and B(7)) xor (A(11) and B(6)) xor (A(12) and B(5)) xor (A(13) and B(4)) xor (A(14) and B(3)) xor (A(15) and B(2)) xor (A(16) and B(1)) xor (A(17) and B(0)) xor (A(10) and B(127)) xor (A(11) and B(126)) xor (A(12) and B(125)) xor (A(13) and B(124)) xor (A(14) and B(123)) xor (A(15) and B(122)) xor (A(16) and B(121)) xor (A(17) and B(120)) xor (A(18) and B(119)) xor (A(19) and B(118)) xor (A(20) and B(117)) xor (A(21) and B(116)) xor (A(23) and B(115)) xor (A(23) and B(114)) xor (A(24) and B(113)) xor (A(25) and B(112)) xor (A(26) and B(111)) xor (A(27) and B(110)) xor (A(28) and B(109)) xor (A(29) and B(108)) xor (A(30) and B(107)) xor (A(31) and B(106)) xor (A(32) and B(105)) xor (A(33) and B(104)) xor (A(34) and B(103)) xor (A(35) and B(102)) xor (A(36) and B(101)) xor (A(37) and B(100)) xor (A(38) and B(99)) xor (A(39) and B(98)) xor (A(40) and B(97)) xor (A(41) and B(96)) xor (A(42) and B(95)) xor (A(43) and B(94)) xor (A(44) and B(93)) xor (A(45) and B(92)) xor (A(46) and B(91)) xor (A(47) and B(90)) xor (A(48) and B(89)) xor (A(49) and B(88)) xor (A(50) and B(87)) xor (A(51) and B(86)) xor (A(52) and B(85)) xor (A(53) and B(84)) xor (A(54) and B(83)) xor (A(55) and B(82)) xor (A(56) and B(81)) xor (A(57) and B(80)) xor (A(58) and B(79)) xor (A(59) and B(78)) xor (A(60) and B(77)) xor (A(61) and B(76)) xor (A(62) and B(75)) xor (A(63) and B(74)) xor (A(64) and B(73)) xor (A(65) and B(72)) xor (A(66) and B(71)) xor (A(67) and B(70)) xor (A(68) and B(69)) xor (A(69) and B(68)) xor (A(70) and B(67)) xor (A(71) and B(66)) xor (A(72) and B(65)) xor (A(73) and B(64)) xor (A(74) and B(63)) xor (A(75) and B(62)) xor (A(76) and B(61)) xor (A(77) and B(60)) xor (A(78) and B(59)) xor (A(79) and B(58)) xor (A(80) and B(57)) xor (A(81) and B(56)) xor (A(82) and B(55)) xor (A(83) and B(54)) xor (A(84) and B(53)) xor (A(85) and B(52)) xor (A(86) and B(51)) xor (A(87) and B(50)) xor (A(88) and B(49)) xor (A(89) and B(48)) xor (A(90) and B(47)) xor (A(91) and B(46)) xor (A(92) and B(45)) xor (A(93) and B(44)) xor (A(94) and B(43)) xor (A(95) and B(42)) xor (A(96) and B(41)) xor (A(97) and B(40)) xor (A(98) and B(39)) xor (A(99) and B(38)) xor (A(100) and B(37)) xor (A(101) and B(36)) xor (A(102) and B(35)) xor (A(103) and B(34)) xor (A(104) and B(33)) xor (A(105) and B(32)) xor (A(106) and B(31)) xor (A(107) and B(30)) xor (A(108) and B(29)) xor (A(109) and B(28)) xor (A(110) and B(27)) xor (A(111) and B(26)) xor (A(112) and B(25)) xor (A(113) and B(24)) xor (A(114) and B(23)) xor (A(115) and B(23)) xor (A(116) and B(21)) xor (A(117) and B(20)) xor (A(118) and B(19)) xor (A(119) and B(18)) xor (A(120) and B(17)) xor (A(121) and B(16)) xor (A(122) and B(15)) xor (A(123) and B(14)) xor (A(124) and B(13)) xor (A(125) and B(12)) xor (A(126) and B(11)) xor (A(15) and B(127)) xor (A(16) and B(126)) xor (A(17) and B(125)) xor (A(18) and B(124)) xor (A(19) and B(123)) xor (A(20) and B(122)) xor (A(21) and B(121)) xor (A(23) and B(120)) xor (A(23) and B(119)) xor (A(24) and B(118)) xor (A(25) and B(117)) xor (A(26) and B(116)) xor (A(27) and B(115)) xor (A(28) and B(114)) xor (A(29) and B(113)) xor (A(30) and B(112)) xor (A(31) and B(111)) xor (A(32) and B(110)) xor (A(33) and B(109)) xor (A(34) and B(108)) xor (A(35) and B(107)) xor (A(36) and B(106)) xor (A(37) and B(105)) xor (A(38) and B(104)) xor (A(39) and B(103)) xor (A(40) and B(102)) xor (A(41) and B(101)) xor (A(42) and B(100)) xor (A(43) and B(99)) xor (A(44) and B(98)) xor (A(45) and B(97)) xor (A(46) and B(96)) xor (A(47) and B(95)) xor (A(48) and B(94)) xor (A(49) and B(93)) xor (A(50) and B(92)) xor (A(51) and B(91)) xor (A(52) and B(90)) xor (A(53) and B(89)) xor (A(54) and B(88)) xor (A(55) and B(87)) xor (A(56) and B(86)) xor (A(57) and B(85)) xor (A(58) and B(84)) xor (A(59) and B(83)) xor (A(60) and B(82)) xor (A(61) and B(81)) xor (A(62) and B(80)) xor (A(63) and B(79)) xor (A(64) and B(78)) xor (A(65) and B(77)) xor (A(66) and B(76)) xor (A(67) and B(75)) xor (A(68) and B(74)) xor (A(69) and B(73)) xor (A(70) and B(72)) xor (A(71) and B(71)) xor (A(72) and B(70)) xor (A(73) and B(69)) xor (A(74) and B(68)) xor (A(75) and B(67)) xor (A(76) and B(66)) xor (A(77) and B(65)) xor (A(78) and B(64)) xor (A(79) and B(63)) xor (A(80) and B(62)) xor (A(81) and B(61)) xor (A(82) and B(60)) xor (A(83) and B(59)) xor (A(84) and B(58)) xor (A(85) and B(57)) xor (A(86) and B(56)) xor (A(87) and B(55)) xor (A(88) and B(54)) xor (A(89) and B(53)) xor (A(90) and B(52)) xor (A(91) and B(51)) xor (A(92) and B(50)) xor (A(93) and B(49)) xor (A(94) and B(48)) xor (A(95) and B(47)) xor (A(96) and B(46)) xor (A(97) and B(45)) xor (A(98) and B(44)) xor (A(99) and B(43)) xor (A(100) and B(42)) xor (A(101) and B(41)) xor (A(102) and B(40)) xor (A(103) and B(39)) xor (A(104) and B(38)) xor (A(105) and B(37)) xor (A(106) and B(36)) xor (A(107) and B(35)) xor (A(108) and B(34)) xor (A(109) and B(33)) xor (A(110) and B(32)) xor (A(111) and B(31)) xor (A(112) and B(30)) xor (A(113) and B(29)) xor (A(114) and B(28)) xor (A(115) and B(27)) xor (A(116) and B(26)) xor (A(117) and B(25)) xor (A(118) and B(24)) xor (A(119) and B(23)) xor (A(120) and B(23)) xor (A(121) and B(21)) xor (A(122) and B(20)) xor (A(123) and B(19)) xor (A(124) and B(18)) xor (A(125) and B(17)) xor (A(126) and B(16)) xor (A(16) and B(127)) xor (A(17) and B(126)) xor (A(18) and B(125)) xor (A(19) and B(124)) xor (A(20) and B(123)) xor (A(21) and B(122)) xor (A(23) and B(121)) xor (A(23) and B(120)) xor (A(24) and B(119)) xor (A(25) and B(118)) xor (A(26) and B(117)) xor (A(27) and B(116)) xor (A(28) and B(115)) xor (A(29) and B(114)) xor (A(30) and B(113)) xor (A(31) and B(112)) xor (A(32) and B(111)) xor (A(33) and B(110)) xor (A(34) and B(109)) xor (A(35) and B(108)) xor (A(36) and B(107)) xor (A(37) and B(106)) xor (A(38) and B(105)) xor (A(39) and B(104)) xor (A(40) and B(103)) xor (A(41) and B(102)) xor (A(42) and B(101)) xor (A(43) and B(100)) xor (A(44) and B(99)) xor (A(45) and B(98)) xor (A(46) and B(97)) xor (A(47) and B(96)) xor (A(48) and B(95)) xor (A(49) and B(94)) xor (A(50) and B(93)) xor (A(51) and B(92)) xor (A(52) and B(91)) xor (A(53) and B(90)) xor (A(54) and B(89)) xor (A(55) and B(88)) xor (A(56) and B(87)) xor (A(57) and B(86)) xor (A(58) and B(85)) xor (A(59) and B(84)) xor (A(60) and B(83)) xor (A(61) and B(82)) xor (A(62) and B(81)) xor (A(63) and B(80)) xor (A(64) and B(79)) xor (A(65) and B(78)) xor (A(66) and B(77)) xor (A(67) and B(76)) xor (A(68) and B(75)) xor (A(69) and B(74)) xor (A(70) and B(73)) xor (A(71) and B(72)) xor (A(72) and B(71)) xor (A(73) and B(70)) xor (A(74) and B(69)) xor (A(75) and B(68)) xor (A(76) and B(67)) xor (A(77) and B(66)) xor (A(78) and B(65)) xor (A(79) and B(64)) xor (A(80) and B(63)) xor (A(81) and B(62)) xor (A(82) and B(61)) xor (A(83) and B(60)) xor (A(84) and B(59)) xor (A(85) and B(58)) xor (A(86) and B(57)) xor (A(87) and B(56)) xor (A(88) and B(55)) xor (A(89) and B(54)) xor (A(90) and B(53)) xor (A(91) and B(52)) xor (A(92) and B(51)) xor (A(93) and B(50)) xor (A(94) and B(49)) xor (A(95) and B(48)) xor (A(96) and B(47)) xor (A(97) and B(46)) xor (A(98) and B(45)) xor (A(99) and B(44)) xor (A(100) and B(43)) xor (A(101) and B(42)) xor (A(102) and B(41)) xor (A(103) and B(40)) xor (A(104) and B(39)) xor (A(105) and B(38)) xor (A(106) and B(37)) xor (A(107) and B(36)) xor (A(108) and B(35)) xor (A(109) and B(34)) xor (A(110) and B(33)) xor (A(111) and B(32)) xor (A(112) and B(31)) xor (A(113) and B(30)) xor (A(114) and B(29)) xor (A(115) and B(28)) xor (A(116) and B(27)) xor (A(117) and B(26)) xor (A(118) and B(25)) xor (A(119) and B(24)) xor (A(120) and B(23)) xor (A(121) and B(23)) xor (A(122) and B(21)) xor (A(123) and B(20)) xor (A(124) and B(19)) xor (A(125) and B(18)) xor (A(126) and B(17)) xor (A(17) and B(127)) xor (A(18) and B(126)) xor (A(19) and B(125)) xor (A(20) and B(124)) xor (A(21) and B(123)) xor (A(23) and B(122)) xor (A(23) and B(121)) xor (A(24) and B(120)) xor (A(25) and B(119)) xor (A(26) and B(118)) xor (A(27) and B(117)) xor (A(28) and B(116)) xor (A(29) and B(115)) xor (A(30) and B(114)) xor (A(31) and B(113)) xor (A(32) and B(112)) xor (A(33) and B(111)) xor (A(34) and B(110)) xor (A(35) and B(109)) xor (A(36) and B(108)) xor (A(37) and B(107)) xor (A(38) and B(106)) xor (A(39) and B(105)) xor (A(40) and B(104)) xor (A(41) and B(103)) xor (A(42) and B(102)) xor (A(43) and B(101)) xor (A(44) and B(100)) xor (A(45) and B(99)) xor (A(46) and B(98)) xor (A(47) and B(97)) xor (A(48) and B(96)) xor (A(49) and B(95)) xor (A(50) and B(94)) xor (A(51) and B(93)) xor (A(52) and B(92)) xor (A(53) and B(91)) xor (A(54) and B(90)) xor (A(55) and B(89)) xor (A(56) and B(88)) xor (A(57) and B(87)) xor (A(58) and B(86)) xor (A(59) and B(85)) xor (A(60) and B(84)) xor (A(61) and B(83)) xor (A(62) and B(82)) xor (A(63) and B(81)) xor (A(64) and B(80)) xor (A(65) and B(79)) xor (A(66) and B(78)) xor (A(67) and B(77)) xor (A(68) and B(76)) xor (A(69) and B(75)) xor (A(70) and B(74)) xor (A(71) and B(73)) xor (A(72) and B(72)) xor (A(73) and B(71)) xor (A(74) and B(70)) xor (A(75) and B(69)) xor (A(76) and B(68)) xor (A(77) and B(67)) xor (A(78) and B(66)) xor (A(79) and B(65)) xor (A(80) and B(64)) xor (A(81) and B(63)) xor (A(82) and B(62)) xor (A(83) and B(61)) xor (A(84) and B(60)) xor (A(85) and B(59)) xor (A(86) and B(58)) xor (A(87) and B(57)) xor (A(88) and B(56)) xor (A(89) and B(55)) xor (A(90) and B(54)) xor (A(91) and B(53)) xor (A(92) and B(52)) xor (A(93) and B(51)) xor (A(94) and B(50)) xor (A(95) and B(49)) xor (A(96) and B(48)) xor (A(97) and B(47)) xor (A(98) and B(46)) xor (A(99) and B(45)) xor (A(100) and B(44)) xor (A(101) and B(43)) xor (A(102) and B(42)) xor (A(103) and B(41)) xor (A(104) and B(40)) xor (A(105) and B(39)) xor (A(106) and B(38)) xor (A(107) and B(37)) xor (A(108) and B(36)) xor (A(109) and B(35)) xor (A(110) and B(34)) xor (A(111) and B(33)) xor (A(112) and B(32)) xor (A(113) and B(31)) xor (A(114) and B(30)) xor (A(115) and B(29)) xor (A(116) and B(28)) xor (A(117) and B(27)) xor (A(118) and B(26)) xor (A(119) and B(25)) xor (A(120) and B(24)) xor (A(121) and B(23)) xor (A(122) and B(23)) xor (A(123) and B(21)) xor (A(124) and B(20)) xor (A(125) and B(19)) xor (A(126) and B(19));
    C(18)  <= (A(0) and B(18)) xor (A(1) and B(17)) xor (A(2) and B(16)) xor (A(3) and B(15)) xor (A(4) and B(14)) xor (A(5) and B(13)) xor (A(6) and B(12)) xor (A(7) and B(11)) xor (A(8) and B(10)) xor (A(9) and B(9)) xor (A(10) and B(8)) xor (A(11) and B(7)) xor (A(12) and B(6)) xor (A(13) and B(5)) xor (A(14) and B(4)) xor (A(15) and B(3)) xor (A(16) and B(2)) xor (A(17) and B(1)) xor (A(18) and B(0)) xor (A(11) and B(127)) xor (A(12) and B(126)) xor (A(13) and B(125)) xor (A(14) and B(124)) xor (A(15) and B(123)) xor (A(16) and B(122)) xor (A(17) and B(121)) xor (A(18) and B(120)) xor (A(19) and B(119)) xor (A(20) and B(118)) xor (A(21) and B(117)) xor (A(23) and B(116)) xor (A(23) and B(115)) xor (A(24) and B(114)) xor (A(25) and B(113)) xor (A(26) and B(112)) xor (A(27) and B(111)) xor (A(28) and B(110)) xor (A(29) and B(109)) xor (A(30) and B(108)) xor (A(31) and B(107)) xor (A(32) and B(106)) xor (A(33) and B(105)) xor (A(34) and B(104)) xor (A(35) and B(103)) xor (A(36) and B(102)) xor (A(37) and B(101)) xor (A(38) and B(100)) xor (A(39) and B(99)) xor (A(40) and B(98)) xor (A(41) and B(97)) xor (A(42) and B(96)) xor (A(43) and B(95)) xor (A(44) and B(94)) xor (A(45) and B(93)) xor (A(46) and B(92)) xor (A(47) and B(91)) xor (A(48) and B(90)) xor (A(49) and B(89)) xor (A(50) and B(88)) xor (A(51) and B(87)) xor (A(52) and B(86)) xor (A(53) and B(85)) xor (A(54) and B(84)) xor (A(55) and B(83)) xor (A(56) and B(82)) xor (A(57) and B(81)) xor (A(58) and B(80)) xor (A(59) and B(79)) xor (A(60) and B(78)) xor (A(61) and B(77)) xor (A(62) and B(76)) xor (A(63) and B(75)) xor (A(64) and B(74)) xor (A(65) and B(73)) xor (A(66) and B(72)) xor (A(67) and B(71)) xor (A(68) and B(70)) xor (A(69) and B(69)) xor (A(70) and B(68)) xor (A(71) and B(67)) xor (A(72) and B(66)) xor (A(73) and B(65)) xor (A(74) and B(64)) xor (A(75) and B(63)) xor (A(76) and B(62)) xor (A(77) and B(61)) xor (A(78) and B(60)) xor (A(79) and B(59)) xor (A(80) and B(58)) xor (A(81) and B(57)) xor (A(82) and B(56)) xor (A(83) and B(55)) xor (A(84) and B(54)) xor (A(85) and B(53)) xor (A(86) and B(52)) xor (A(87) and B(51)) xor (A(88) and B(50)) xor (A(89) and B(49)) xor (A(90) and B(48)) xor (A(91) and B(47)) xor (A(92) and B(46)) xor (A(93) and B(45)) xor (A(94) and B(44)) xor (A(95) and B(43)) xor (A(96) and B(42)) xor (A(97) and B(41)) xor (A(98) and B(40)) xor (A(99) and B(39)) xor (A(100) and B(38)) xor (A(101) and B(37)) xor (A(102) and B(36)) xor (A(103) and B(35)) xor (A(104) and B(34)) xor (A(105) and B(33)) xor (A(106) and B(32)) xor (A(107) and B(31)) xor (A(108) and B(30)) xor (A(109) and B(29)) xor (A(110) and B(28)) xor (A(111) and B(27)) xor (A(112) and B(26)) xor (A(113) and B(25)) xor (A(114) and B(24)) xor (A(115) and B(23)) xor (A(116) and B(23)) xor (A(117) and B(21)) xor (A(118) and B(20)) xor (A(119) and B(19)) xor (A(120) and B(18)) xor (A(121) and B(17)) xor (A(122) and B(16)) xor (A(123) and B(15)) xor (A(124) and B(14)) xor (A(125) and B(13)) xor (A(126) and B(12)) xor (A(16) and B(127)) xor (A(17) and B(126)) xor (A(18) and B(125)) xor (A(19) and B(124)) xor (A(20) and B(123)) xor (A(21) and B(122)) xor (A(23) and B(121)) xor (A(23) and B(120)) xor (A(24) and B(119)) xor (A(25) and B(118)) xor (A(26) and B(117)) xor (A(27) and B(116)) xor (A(28) and B(115)) xor (A(29) and B(114)) xor (A(30) and B(113)) xor (A(31) and B(112)) xor (A(32) and B(111)) xor (A(33) and B(110)) xor (A(34) and B(109)) xor (A(35) and B(108)) xor (A(36) and B(107)) xor (A(37) and B(106)) xor (A(38) and B(105)) xor (A(39) and B(104)) xor (A(40) and B(103)) xor (A(41) and B(102)) xor (A(42) and B(101)) xor (A(43) and B(100)) xor (A(44) and B(99)) xor (A(45) and B(98)) xor (A(46) and B(97)) xor (A(47) and B(96)) xor (A(48) and B(95)) xor (A(49) and B(94)) xor (A(50) and B(93)) xor (A(51) and B(92)) xor (A(52) and B(91)) xor (A(53) and B(90)) xor (A(54) and B(89)) xor (A(55) and B(88)) xor (A(56) and B(87)) xor (A(57) and B(86)) xor (A(58) and B(85)) xor (A(59) and B(84)) xor (A(60) and B(83)) xor (A(61) and B(82)) xor (A(62) and B(81)) xor (A(63) and B(80)) xor (A(64) and B(79)) xor (A(65) and B(78)) xor (A(66) and B(77)) xor (A(67) and B(76)) xor (A(68) and B(75)) xor (A(69) and B(74)) xor (A(70) and B(73)) xor (A(71) and B(72)) xor (A(72) and B(71)) xor (A(73) and B(70)) xor (A(74) and B(69)) xor (A(75) and B(68)) xor (A(76) and B(67)) xor (A(77) and B(66)) xor (A(78) and B(65)) xor (A(79) and B(64)) xor (A(80) and B(63)) xor (A(81) and B(62)) xor (A(82) and B(61)) xor (A(83) and B(60)) xor (A(84) and B(59)) xor (A(85) and B(58)) xor (A(86) and B(57)) xor (A(87) and B(56)) xor (A(88) and B(55)) xor (A(89) and B(54)) xor (A(90) and B(53)) xor (A(91) and B(52)) xor (A(92) and B(51)) xor (A(93) and B(50)) xor (A(94) and B(49)) xor (A(95) and B(48)) xor (A(96) and B(47)) xor (A(97) and B(46)) xor (A(98) and B(45)) xor (A(99) and B(44)) xor (A(100) and B(43)) xor (A(101) and B(42)) xor (A(102) and B(41)) xor (A(103) and B(40)) xor (A(104) and B(39)) xor (A(105) and B(38)) xor (A(106) and B(37)) xor (A(107) and B(36)) xor (A(108) and B(35)) xor (A(109) and B(34)) xor (A(110) and B(33)) xor (A(111) and B(32)) xor (A(112) and B(31)) xor (A(113) and B(30)) xor (A(114) and B(29)) xor (A(115) and B(28)) xor (A(116) and B(27)) xor (A(117) and B(26)) xor (A(118) and B(25)) xor (A(119) and B(24)) xor (A(120) and B(23)) xor (A(121) and B(23)) xor (A(122) and B(21)) xor (A(123) and B(20)) xor (A(124) and B(19)) xor (A(125) and B(18)) xor (A(126) and B(17)) xor (A(17) and B(127)) xor (A(18) and B(126)) xor (A(19) and B(125)) xor (A(20) and B(124)) xor (A(21) and B(123)) xor (A(23) and B(122)) xor (A(23) and B(121)) xor (A(24) and B(120)) xor (A(25) and B(119)) xor (A(26) and B(118)) xor (A(27) and B(117)) xor (A(28) and B(116)) xor (A(29) and B(115)) xor (A(30) and B(114)) xor (A(31) and B(113)) xor (A(32) and B(112)) xor (A(33) and B(111)) xor (A(34) and B(110)) xor (A(35) and B(109)) xor (A(36) and B(108)) xor (A(37) and B(107)) xor (A(38) and B(106)) xor (A(39) and B(105)) xor (A(40) and B(104)) xor (A(41) and B(103)) xor (A(42) and B(102)) xor (A(43) and B(101)) xor (A(44) and B(100)) xor (A(45) and B(99)) xor (A(46) and B(98)) xor (A(47) and B(97)) xor (A(48) and B(96)) xor (A(49) and B(95)) xor (A(50) and B(94)) xor (A(51) and B(93)) xor (A(52) and B(92)) xor (A(53) and B(91)) xor (A(54) and B(90)) xor (A(55) and B(89)) xor (A(56) and B(88)) xor (A(57) and B(87)) xor (A(58) and B(86)) xor (A(59) and B(85)) xor (A(60) and B(84)) xor (A(61) and B(83)) xor (A(62) and B(82)) xor (A(63) and B(81)) xor (A(64) and B(80)) xor (A(65) and B(79)) xor (A(66) and B(78)) xor (A(67) and B(77)) xor (A(68) and B(76)) xor (A(69) and B(75)) xor (A(70) and B(74)) xor (A(71) and B(73)) xor (A(72) and B(72)) xor (A(73) and B(71)) xor (A(74) and B(70)) xor (A(75) and B(69)) xor (A(76) and B(68)) xor (A(77) and B(67)) xor (A(78) and B(66)) xor (A(79) and B(65)) xor (A(80) and B(64)) xor (A(81) and B(63)) xor (A(82) and B(62)) xor (A(83) and B(61)) xor (A(84) and B(60)) xor (A(85) and B(59)) xor (A(86) and B(58)) xor (A(87) and B(57)) xor (A(88) and B(56)) xor (A(89) and B(55)) xor (A(90) and B(54)) xor (A(91) and B(53)) xor (A(92) and B(52)) xor (A(93) and B(51)) xor (A(94) and B(50)) xor (A(95) and B(49)) xor (A(96) and B(48)) xor (A(97) and B(47)) xor (A(98) and B(46)) xor (A(99) and B(45)) xor (A(100) and B(44)) xor (A(101) and B(43)) xor (A(102) and B(42)) xor (A(103) and B(41)) xor (A(104) and B(40)) xor (A(105) and B(39)) xor (A(106) and B(38)) xor (A(107) and B(37)) xor (A(108) and B(36)) xor (A(109) and B(35)) xor (A(110) and B(34)) xor (A(111) and B(33)) xor (A(112) and B(32)) xor (A(113) and B(31)) xor (A(114) and B(30)) xor (A(115) and B(29)) xor (A(116) and B(28)) xor (A(117) and B(27)) xor (A(118) and B(26)) xor (A(119) and B(25)) xor (A(120) and B(24)) xor (A(121) and B(23)) xor (A(122) and B(23)) xor (A(123) and B(21)) xor (A(124) and B(20)) xor (A(125) and B(19)) xor (A(126) and B(18)) xor (A(18) and B(127)) xor (A(19) and B(126)) xor (A(20) and B(125)) xor (A(21) and B(124)) xor (A(23) and B(123)) xor (A(23) and B(122)) xor (A(24) and B(121)) xor (A(25) and B(120)) xor (A(26) and B(119)) xor (A(27) and B(118)) xor (A(28) and B(117)) xor (A(29) and B(116)) xor (A(30) and B(115)) xor (A(31) and B(114)) xor (A(32) and B(113)) xor (A(33) and B(112)) xor (A(34) and B(111)) xor (A(35) and B(110)) xor (A(36) and B(109)) xor (A(37) and B(108)) xor (A(38) and B(107)) xor (A(39) and B(106)) xor (A(40) and B(105)) xor (A(41) and B(104)) xor (A(42) and B(103)) xor (A(43) and B(102)) xor (A(44) and B(101)) xor (A(45) and B(100)) xor (A(46) and B(99)) xor (A(47) and B(98)) xor (A(48) and B(97)) xor (A(49) and B(96)) xor (A(50) and B(95)) xor (A(51) and B(94)) xor (A(52) and B(93)) xor (A(53) and B(92)) xor (A(54) and B(91)) xor (A(55) and B(90)) xor (A(56) and B(89)) xor (A(57) and B(88)) xor (A(58) and B(87)) xor (A(59) and B(86)) xor (A(60) and B(85)) xor (A(61) and B(84)) xor (A(62) and B(83)) xor (A(63) and B(82)) xor (A(64) and B(81)) xor (A(65) and B(80)) xor (A(66) and B(79)) xor (A(67) and B(78)) xor (A(68) and B(77)) xor (A(69) and B(76)) xor (A(70) and B(75)) xor (A(71) and B(74)) xor (A(72) and B(73)) xor (A(73) and B(72)) xor (A(74) and B(71)) xor (A(75) and B(70)) xor (A(76) and B(69)) xor (A(77) and B(68)) xor (A(78) and B(67)) xor (A(79) and B(66)) xor (A(80) and B(65)) xor (A(81) and B(64)) xor (A(82) and B(63)) xor (A(83) and B(62)) xor (A(84) and B(61)) xor (A(85) and B(60)) xor (A(86) and B(59)) xor (A(87) and B(58)) xor (A(88) and B(57)) xor (A(89) and B(56)) xor (A(90) and B(55)) xor (A(91) and B(54)) xor (A(92) and B(53)) xor (A(93) and B(52)) xor (A(94) and B(51)) xor (A(95) and B(50)) xor (A(96) and B(49)) xor (A(97) and B(48)) xor (A(98) and B(47)) xor (A(99) and B(46)) xor (A(100) and B(45)) xor (A(101) and B(44)) xor (A(102) and B(43)) xor (A(103) and B(42)) xor (A(104) and B(41)) xor (A(105) and B(40)) xor (A(106) and B(39)) xor (A(107) and B(38)) xor (A(108) and B(37)) xor (A(109) and B(36)) xor (A(110) and B(35)) xor (A(111) and B(34)) xor (A(112) and B(33)) xor (A(113) and B(32)) xor (A(114) and B(31)) xor (A(115) and B(30)) xor (A(116) and B(29)) xor (A(117) and B(28)) xor (A(118) and B(27)) xor (A(119) and B(26)) xor (A(120) and B(25)) xor (A(121) and B(24)) xor (A(122) and B(23)) xor (A(123) and B(23)) xor (A(124) and B(21)) xor (A(125) and B(20)) xor (A(126) and B(20));
    C(19)  <= (A(0) and B(19)) xor (A(1) and B(18)) xor (A(2) and B(17)) xor (A(3) and B(16)) xor (A(4) and B(15)) xor (A(5) and B(14)) xor (A(6) and B(13)) xor (A(7) and B(12)) xor (A(8) and B(11)) xor (A(9) and B(10)) xor (A(10) and B(9)) xor (A(11) and B(8)) xor (A(12) and B(7)) xor (A(13) and B(6)) xor (A(14) and B(5)) xor (A(15) and B(4)) xor (A(16) and B(3)) xor (A(17) and B(2)) xor (A(18) and B(1)) xor (A(19) and B(0)) xor (A(12) and B(127)) xor (A(13) and B(126)) xor (A(14) and B(125)) xor (A(15) and B(124)) xor (A(16) and B(123)) xor (A(17) and B(122)) xor (A(18) and B(121)) xor (A(19) and B(120)) xor (A(20) and B(119)) xor (A(21) and B(118)) xor (A(23) and B(117)) xor (A(23) and B(116)) xor (A(24) and B(115)) xor (A(25) and B(114)) xor (A(26) and B(113)) xor (A(27) and B(112)) xor (A(28) and B(111)) xor (A(29) and B(110)) xor (A(30) and B(109)) xor (A(31) and B(108)) xor (A(32) and B(107)) xor (A(33) and B(106)) xor (A(34) and B(105)) xor (A(35) and B(104)) xor (A(36) and B(103)) xor (A(37) and B(102)) xor (A(38) and B(101)) xor (A(39) and B(100)) xor (A(40) and B(99)) xor (A(41) and B(98)) xor (A(42) and B(97)) xor (A(43) and B(96)) xor (A(44) and B(95)) xor (A(45) and B(94)) xor (A(46) and B(93)) xor (A(47) and B(92)) xor (A(48) and B(91)) xor (A(49) and B(90)) xor (A(50) and B(89)) xor (A(51) and B(88)) xor (A(52) and B(87)) xor (A(53) and B(86)) xor (A(54) and B(85)) xor (A(55) and B(84)) xor (A(56) and B(83)) xor (A(57) and B(82)) xor (A(58) and B(81)) xor (A(59) and B(80)) xor (A(60) and B(79)) xor (A(61) and B(78)) xor (A(62) and B(77)) xor (A(63) and B(76)) xor (A(64) and B(75)) xor (A(65) and B(74)) xor (A(66) and B(73)) xor (A(67) and B(72)) xor (A(68) and B(71)) xor (A(69) and B(70)) xor (A(70) and B(69)) xor (A(71) and B(68)) xor (A(72) and B(67)) xor (A(73) and B(66)) xor (A(74) and B(65)) xor (A(75) and B(64)) xor (A(76) and B(63)) xor (A(77) and B(62)) xor (A(78) and B(61)) xor (A(79) and B(60)) xor (A(80) and B(59)) xor (A(81) and B(58)) xor (A(82) and B(57)) xor (A(83) and B(56)) xor (A(84) and B(55)) xor (A(85) and B(54)) xor (A(86) and B(53)) xor (A(87) and B(52)) xor (A(88) and B(51)) xor (A(89) and B(50)) xor (A(90) and B(49)) xor (A(91) and B(48)) xor (A(92) and B(47)) xor (A(93) and B(46)) xor (A(94) and B(45)) xor (A(95) and B(44)) xor (A(96) and B(43)) xor (A(97) and B(42)) xor (A(98) and B(41)) xor (A(99) and B(40)) xor (A(100) and B(39)) xor (A(101) and B(38)) xor (A(102) and B(37)) xor (A(103) and B(36)) xor (A(104) and B(35)) xor (A(105) and B(34)) xor (A(106) and B(33)) xor (A(107) and B(32)) xor (A(108) and B(31)) xor (A(109) and B(30)) xor (A(110) and B(29)) xor (A(111) and B(28)) xor (A(112) and B(27)) xor (A(113) and B(26)) xor (A(114) and B(25)) xor (A(115) and B(24)) xor (A(116) and B(23)) xor (A(117) and B(23)) xor (A(118) and B(21)) xor (A(119) and B(20)) xor (A(120) and B(19)) xor (A(121) and B(18)) xor (A(122) and B(17)) xor (A(123) and B(16)) xor (A(124) and B(15)) xor (A(125) and B(14)) xor (A(126) and B(13)) xor (A(17) and B(127)) xor (A(18) and B(126)) xor (A(19) and B(125)) xor (A(20) and B(124)) xor (A(21) and B(123)) xor (A(23) and B(122)) xor (A(23) and B(121)) xor (A(24) and B(120)) xor (A(25) and B(119)) xor (A(26) and B(118)) xor (A(27) and B(117)) xor (A(28) and B(116)) xor (A(29) and B(115)) xor (A(30) and B(114)) xor (A(31) and B(113)) xor (A(32) and B(112)) xor (A(33) and B(111)) xor (A(34) and B(110)) xor (A(35) and B(109)) xor (A(36) and B(108)) xor (A(37) and B(107)) xor (A(38) and B(106)) xor (A(39) and B(105)) xor (A(40) and B(104)) xor (A(41) and B(103)) xor (A(42) and B(102)) xor (A(43) and B(101)) xor (A(44) and B(100)) xor (A(45) and B(99)) xor (A(46) and B(98)) xor (A(47) and B(97)) xor (A(48) and B(96)) xor (A(49) and B(95)) xor (A(50) and B(94)) xor (A(51) and B(93)) xor (A(52) and B(92)) xor (A(53) and B(91)) xor (A(54) and B(90)) xor (A(55) and B(89)) xor (A(56) and B(88)) xor (A(57) and B(87)) xor (A(58) and B(86)) xor (A(59) and B(85)) xor (A(60) and B(84)) xor (A(61) and B(83)) xor (A(62) and B(82)) xor (A(63) and B(81)) xor (A(64) and B(80)) xor (A(65) and B(79)) xor (A(66) and B(78)) xor (A(67) and B(77)) xor (A(68) and B(76)) xor (A(69) and B(75)) xor (A(70) and B(74)) xor (A(71) and B(73)) xor (A(72) and B(72)) xor (A(73) and B(71)) xor (A(74) and B(70)) xor (A(75) and B(69)) xor (A(76) and B(68)) xor (A(77) and B(67)) xor (A(78) and B(66)) xor (A(79) and B(65)) xor (A(80) and B(64)) xor (A(81) and B(63)) xor (A(82) and B(62)) xor (A(83) and B(61)) xor (A(84) and B(60)) xor (A(85) and B(59)) xor (A(86) and B(58)) xor (A(87) and B(57)) xor (A(88) and B(56)) xor (A(89) and B(55)) xor (A(90) and B(54)) xor (A(91) and B(53)) xor (A(92) and B(52)) xor (A(93) and B(51)) xor (A(94) and B(50)) xor (A(95) and B(49)) xor (A(96) and B(48)) xor (A(97) and B(47)) xor (A(98) and B(46)) xor (A(99) and B(45)) xor (A(100) and B(44)) xor (A(101) and B(43)) xor (A(102) and B(42)) xor (A(103) and B(41)) xor (A(104) and B(40)) xor (A(105) and B(39)) xor (A(106) and B(38)) xor (A(107) and B(37)) xor (A(108) and B(36)) xor (A(109) and B(35)) xor (A(110) and B(34)) xor (A(111) and B(33)) xor (A(112) and B(32)) xor (A(113) and B(31)) xor (A(114) and B(30)) xor (A(115) and B(29)) xor (A(116) and B(28)) xor (A(117) and B(27)) xor (A(118) and B(26)) xor (A(119) and B(25)) xor (A(120) and B(24)) xor (A(121) and B(23)) xor (A(122) and B(23)) xor (A(123) and B(21)) xor (A(124) and B(20)) xor (A(125) and B(19)) xor (A(126) and B(18)) xor (A(18) and B(127)) xor (A(19) and B(126)) xor (A(20) and B(125)) xor (A(21) and B(124)) xor (A(23) and B(123)) xor (A(23) and B(122)) xor (A(24) and B(121)) xor (A(25) and B(120)) xor (A(26) and B(119)) xor (A(27) and B(118)) xor (A(28) and B(117)) xor (A(29) and B(116)) xor (A(30) and B(115)) xor (A(31) and B(114)) xor (A(32) and B(113)) xor (A(33) and B(112)) xor (A(34) and B(111)) xor (A(35) and B(110)) xor (A(36) and B(109)) xor (A(37) and B(108)) xor (A(38) and B(107)) xor (A(39) and B(106)) xor (A(40) and B(105)) xor (A(41) and B(104)) xor (A(42) and B(103)) xor (A(43) and B(102)) xor (A(44) and B(101)) xor (A(45) and B(100)) xor (A(46) and B(99)) xor (A(47) and B(98)) xor (A(48) and B(97)) xor (A(49) and B(96)) xor (A(50) and B(95)) xor (A(51) and B(94)) xor (A(52) and B(93)) xor (A(53) and B(92)) xor (A(54) and B(91)) xor (A(55) and B(90)) xor (A(56) and B(89)) xor (A(57) and B(88)) xor (A(58) and B(87)) xor (A(59) and B(86)) xor (A(60) and B(85)) xor (A(61) and B(84)) xor (A(62) and B(83)) xor (A(63) and B(82)) xor (A(64) and B(81)) xor (A(65) and B(80)) xor (A(66) and B(79)) xor (A(67) and B(78)) xor (A(68) and B(77)) xor (A(69) and B(76)) xor (A(70) and B(75)) xor (A(71) and B(74)) xor (A(72) and B(73)) xor (A(73) and B(72)) xor (A(74) and B(71)) xor (A(75) and B(70)) xor (A(76) and B(69)) xor (A(77) and B(68)) xor (A(78) and B(67)) xor (A(79) and B(66)) xor (A(80) and B(65)) xor (A(81) and B(64)) xor (A(82) and B(63)) xor (A(83) and B(62)) xor (A(84) and B(61)) xor (A(85) and B(60)) xor (A(86) and B(59)) xor (A(87) and B(58)) xor (A(88) and B(57)) xor (A(89) and B(56)) xor (A(90) and B(55)) xor (A(91) and B(54)) xor (A(92) and B(53)) xor (A(93) and B(52)) xor (A(94) and B(51)) xor (A(95) and B(50)) xor (A(96) and B(49)) xor (A(97) and B(48)) xor (A(98) and B(47)) xor (A(99) and B(46)) xor (A(100) and B(45)) xor (A(101) and B(44)) xor (A(102) and B(43)) xor (A(103) and B(42)) xor (A(104) and B(41)) xor (A(105) and B(40)) xor (A(106) and B(39)) xor (A(107) and B(38)) xor (A(108) and B(37)) xor (A(109) and B(36)) xor (A(110) and B(35)) xor (A(111) and B(34)) xor (A(112) and B(33)) xor (A(113) and B(32)) xor (A(114) and B(31)) xor (A(115) and B(30)) xor (A(116) and B(29)) xor (A(117) and B(28)) xor (A(118) and B(27)) xor (A(119) and B(26)) xor (A(120) and B(25)) xor (A(121) and B(24)) xor (A(122) and B(23)) xor (A(123) and B(23)) xor (A(124) and B(21)) xor (A(125) and B(20)) xor (A(126) and B(19)) xor (A(19) and B(127)) xor (A(20) and B(126)) xor (A(21) and B(125)) xor (A(23) and B(124)) xor (A(23) and B(123)) xor (A(24) and B(122)) xor (A(25) and B(121)) xor (A(26) and B(120)) xor (A(27) and B(119)) xor (A(28) and B(118)) xor (A(29) and B(117)) xor (A(30) and B(116)) xor (A(31) and B(115)) xor (A(32) and B(114)) xor (A(33) and B(113)) xor (A(34) and B(112)) xor (A(35) and B(111)) xor (A(36) and B(110)) xor (A(37) and B(109)) xor (A(38) and B(108)) xor (A(39) and B(107)) xor (A(40) and B(106)) xor (A(41) and B(105)) xor (A(42) and B(104)) xor (A(43) and B(103)) xor (A(44) and B(102)) xor (A(45) and B(101)) xor (A(46) and B(100)) xor (A(47) and B(99)) xor (A(48) and B(98)) xor (A(49) and B(97)) xor (A(50) and B(96)) xor (A(51) and B(95)) xor (A(52) and B(94)) xor (A(53) and B(93)) xor (A(54) and B(92)) xor (A(55) and B(91)) xor (A(56) and B(90)) xor (A(57) and B(89)) xor (A(58) and B(88)) xor (A(59) and B(87)) xor (A(60) and B(86)) xor (A(61) and B(85)) xor (A(62) and B(84)) xor (A(63) and B(83)) xor (A(64) and B(82)) xor (A(65) and B(81)) xor (A(66) and B(80)) xor (A(67) and B(79)) xor (A(68) and B(78)) xor (A(69) and B(77)) xor (A(70) and B(76)) xor (A(71) and B(75)) xor (A(72) and B(74)) xor (A(73) and B(73)) xor (A(74) and B(72)) xor (A(75) and B(71)) xor (A(76) and B(70)) xor (A(77) and B(69)) xor (A(78) and B(68)) xor (A(79) and B(67)) xor (A(80) and B(66)) xor (A(81) and B(65)) xor (A(82) and B(64)) xor (A(83) and B(63)) xor (A(84) and B(62)) xor (A(85) and B(61)) xor (A(86) and B(60)) xor (A(87) and B(59)) xor (A(88) and B(58)) xor (A(89) and B(57)) xor (A(90) and B(56)) xor (A(91) and B(55)) xor (A(92) and B(54)) xor (A(93) and B(53)) xor (A(94) and B(52)) xor (A(95) and B(51)) xor (A(96) and B(50)) xor (A(97) and B(49)) xor (A(98) and B(48)) xor (A(99) and B(47)) xor (A(100) and B(46)) xor (A(101) and B(45)) xor (A(102) and B(44)) xor (A(103) and B(43)) xor (A(104) and B(42)) xor (A(105) and B(41)) xor (A(106) and B(40)) xor (A(107) and B(39)) xor (A(108) and B(38)) xor (A(109) and B(37)) xor (A(110) and B(36)) xor (A(111) and B(35)) xor (A(112) and B(34)) xor (A(113) and B(33)) xor (A(114) and B(32)) xor (A(115) and B(31)) xor (A(116) and B(30)) xor (A(117) and B(29)) xor (A(118) and B(28)) xor (A(119) and B(27)) xor (A(120) and B(26)) xor (A(121) and B(25)) xor (A(122) and B(24)) xor (A(123) and B(23)) xor (A(124) and B(23)) xor (A(125) and B(21)) xor (A(126) and B(21));
    C(20)  <= (A(0) and B(20)) xor (A(1) and B(19)) xor (A(2) and B(18)) xor (A(3) and B(17)) xor (A(4) and B(16)) xor (A(5) and B(15)) xor (A(6) and B(14)) xor (A(7) and B(13)) xor (A(8) and B(12)) xor (A(9) and B(11)) xor (A(10) and B(10)) xor (A(11) and B(9)) xor (A(12) and B(8)) xor (A(13) and B(7)) xor (A(14) and B(6)) xor (A(15) and B(5)) xor (A(16) and B(4)) xor (A(17) and B(3)) xor (A(18) and B(2)) xor (A(19) and B(1)) xor (A(20) and B(0)) xor (A(13) and B(127)) xor (A(14) and B(126)) xor (A(15) and B(125)) xor (A(16) and B(124)) xor (A(17) and B(123)) xor (A(18) and B(122)) xor (A(19) and B(121)) xor (A(20) and B(120)) xor (A(21) and B(119)) xor (A(23) and B(118)) xor (A(23) and B(117)) xor (A(24) and B(116)) xor (A(25) and B(115)) xor (A(26) and B(114)) xor (A(27) and B(113)) xor (A(28) and B(112)) xor (A(29) and B(111)) xor (A(30) and B(110)) xor (A(31) and B(109)) xor (A(32) and B(108)) xor (A(33) and B(107)) xor (A(34) and B(106)) xor (A(35) and B(105)) xor (A(36) and B(104)) xor (A(37) and B(103)) xor (A(38) and B(102)) xor (A(39) and B(101)) xor (A(40) and B(100)) xor (A(41) and B(99)) xor (A(42) and B(98)) xor (A(43) and B(97)) xor (A(44) and B(96)) xor (A(45) and B(95)) xor (A(46) and B(94)) xor (A(47) and B(93)) xor (A(48) and B(92)) xor (A(49) and B(91)) xor (A(50) and B(90)) xor (A(51) and B(89)) xor (A(52) and B(88)) xor (A(53) and B(87)) xor (A(54) and B(86)) xor (A(55) and B(85)) xor (A(56) and B(84)) xor (A(57) and B(83)) xor (A(58) and B(82)) xor (A(59) and B(81)) xor (A(60) and B(80)) xor (A(61) and B(79)) xor (A(62) and B(78)) xor (A(63) and B(77)) xor (A(64) and B(76)) xor (A(65) and B(75)) xor (A(66) and B(74)) xor (A(67) and B(73)) xor (A(68) and B(72)) xor (A(69) and B(71)) xor (A(70) and B(70)) xor (A(71) and B(69)) xor (A(72) and B(68)) xor (A(73) and B(67)) xor (A(74) and B(66)) xor (A(75) and B(65)) xor (A(76) and B(64)) xor (A(77) and B(63)) xor (A(78) and B(62)) xor (A(79) and B(61)) xor (A(80) and B(60)) xor (A(81) and B(59)) xor (A(82) and B(58)) xor (A(83) and B(57)) xor (A(84) and B(56)) xor (A(85) and B(55)) xor (A(86) and B(54)) xor (A(87) and B(53)) xor (A(88) and B(52)) xor (A(89) and B(51)) xor (A(90) and B(50)) xor (A(91) and B(49)) xor (A(92) and B(48)) xor (A(93) and B(47)) xor (A(94) and B(46)) xor (A(95) and B(45)) xor (A(96) and B(44)) xor (A(97) and B(43)) xor (A(98) and B(42)) xor (A(99) and B(41)) xor (A(100) and B(40)) xor (A(101) and B(39)) xor (A(102) and B(38)) xor (A(103) and B(37)) xor (A(104) and B(36)) xor (A(105) and B(35)) xor (A(106) and B(34)) xor (A(107) and B(33)) xor (A(108) and B(32)) xor (A(109) and B(31)) xor (A(110) and B(30)) xor (A(111) and B(29)) xor (A(112) and B(28)) xor (A(113) and B(27)) xor (A(114) and B(26)) xor (A(115) and B(25)) xor (A(116) and B(24)) xor (A(117) and B(23)) xor (A(118) and B(23)) xor (A(119) and B(21)) xor (A(120) and B(20)) xor (A(121) and B(19)) xor (A(122) and B(18)) xor (A(123) and B(17)) xor (A(124) and B(16)) xor (A(125) and B(15)) xor (A(126) and B(14)) xor (A(18) and B(127)) xor (A(19) and B(126)) xor (A(20) and B(125)) xor (A(21) and B(124)) xor (A(23) and B(123)) xor (A(23) and B(122)) xor (A(24) and B(121)) xor (A(25) and B(120)) xor (A(26) and B(119)) xor (A(27) and B(118)) xor (A(28) and B(117)) xor (A(29) and B(116)) xor (A(30) and B(115)) xor (A(31) and B(114)) xor (A(32) and B(113)) xor (A(33) and B(112)) xor (A(34) and B(111)) xor (A(35) and B(110)) xor (A(36) and B(109)) xor (A(37) and B(108)) xor (A(38) and B(107)) xor (A(39) and B(106)) xor (A(40) and B(105)) xor (A(41) and B(104)) xor (A(42) and B(103)) xor (A(43) and B(102)) xor (A(44) and B(101)) xor (A(45) and B(100)) xor (A(46) and B(99)) xor (A(47) and B(98)) xor (A(48) and B(97)) xor (A(49) and B(96)) xor (A(50) and B(95)) xor (A(51) and B(94)) xor (A(52) and B(93)) xor (A(53) and B(92)) xor (A(54) and B(91)) xor (A(55) and B(90)) xor (A(56) and B(89)) xor (A(57) and B(88)) xor (A(58) and B(87)) xor (A(59) and B(86)) xor (A(60) and B(85)) xor (A(61) and B(84)) xor (A(62) and B(83)) xor (A(63) and B(82)) xor (A(64) and B(81)) xor (A(65) and B(80)) xor (A(66) and B(79)) xor (A(67) and B(78)) xor (A(68) and B(77)) xor (A(69) and B(76)) xor (A(70) and B(75)) xor (A(71) and B(74)) xor (A(72) and B(73)) xor (A(73) and B(72)) xor (A(74) and B(71)) xor (A(75) and B(70)) xor (A(76) and B(69)) xor (A(77) and B(68)) xor (A(78) and B(67)) xor (A(79) and B(66)) xor (A(80) and B(65)) xor (A(81) and B(64)) xor (A(82) and B(63)) xor (A(83) and B(62)) xor (A(84) and B(61)) xor (A(85) and B(60)) xor (A(86) and B(59)) xor (A(87) and B(58)) xor (A(88) and B(57)) xor (A(89) and B(56)) xor (A(90) and B(55)) xor (A(91) and B(54)) xor (A(92) and B(53)) xor (A(93) and B(52)) xor (A(94) and B(51)) xor (A(95) and B(50)) xor (A(96) and B(49)) xor (A(97) and B(48)) xor (A(98) and B(47)) xor (A(99) and B(46)) xor (A(100) and B(45)) xor (A(101) and B(44)) xor (A(102) and B(43)) xor (A(103) and B(42)) xor (A(104) and B(41)) xor (A(105) and B(40)) xor (A(106) and B(39)) xor (A(107) and B(38)) xor (A(108) and B(37)) xor (A(109) and B(36)) xor (A(110) and B(35)) xor (A(111) and B(34)) xor (A(112) and B(33)) xor (A(113) and B(32)) xor (A(114) and B(31)) xor (A(115) and B(30)) xor (A(116) and B(29)) xor (A(117) and B(28)) xor (A(118) and B(27)) xor (A(119) and B(26)) xor (A(120) and B(25)) xor (A(121) and B(24)) xor (A(122) and B(23)) xor (A(123) and B(23)) xor (A(124) and B(21)) xor (A(125) and B(20)) xor (A(126) and B(19)) xor (A(19) and B(127)) xor (A(20) and B(126)) xor (A(21) and B(125)) xor (A(23) and B(124)) xor (A(23) and B(123)) xor (A(24) and B(122)) xor (A(25) and B(121)) xor (A(26) and B(120)) xor (A(27) and B(119)) xor (A(28) and B(118)) xor (A(29) and B(117)) xor (A(30) and B(116)) xor (A(31) and B(115)) xor (A(32) and B(114)) xor (A(33) and B(113)) xor (A(34) and B(112)) xor (A(35) and B(111)) xor (A(36) and B(110)) xor (A(37) and B(109)) xor (A(38) and B(108)) xor (A(39) and B(107)) xor (A(40) and B(106)) xor (A(41) and B(105)) xor (A(42) and B(104)) xor (A(43) and B(103)) xor (A(44) and B(102)) xor (A(45) and B(101)) xor (A(46) and B(100)) xor (A(47) and B(99)) xor (A(48) and B(98)) xor (A(49) and B(97)) xor (A(50) and B(96)) xor (A(51) and B(95)) xor (A(52) and B(94)) xor (A(53) and B(93)) xor (A(54) and B(92)) xor (A(55) and B(91)) xor (A(56) and B(90)) xor (A(57) and B(89)) xor (A(58) and B(88)) xor (A(59) and B(87)) xor (A(60) and B(86)) xor (A(61) and B(85)) xor (A(62) and B(84)) xor (A(63) and B(83)) xor (A(64) and B(82)) xor (A(65) and B(81)) xor (A(66) and B(80)) xor (A(67) and B(79)) xor (A(68) and B(78)) xor (A(69) and B(77)) xor (A(70) and B(76)) xor (A(71) and B(75)) xor (A(72) and B(74)) xor (A(73) and B(73)) xor (A(74) and B(72)) xor (A(75) and B(71)) xor (A(76) and B(70)) xor (A(77) and B(69)) xor (A(78) and B(68)) xor (A(79) and B(67)) xor (A(80) and B(66)) xor (A(81) and B(65)) xor (A(82) and B(64)) xor (A(83) and B(63)) xor (A(84) and B(62)) xor (A(85) and B(61)) xor (A(86) and B(60)) xor (A(87) and B(59)) xor (A(88) and B(58)) xor (A(89) and B(57)) xor (A(90) and B(56)) xor (A(91) and B(55)) xor (A(92) and B(54)) xor (A(93) and B(53)) xor (A(94) and B(52)) xor (A(95) and B(51)) xor (A(96) and B(50)) xor (A(97) and B(49)) xor (A(98) and B(48)) xor (A(99) and B(47)) xor (A(100) and B(46)) xor (A(101) and B(45)) xor (A(102) and B(44)) xor (A(103) and B(43)) xor (A(104) and B(42)) xor (A(105) and B(41)) xor (A(106) and B(40)) xor (A(107) and B(39)) xor (A(108) and B(38)) xor (A(109) and B(37)) xor (A(110) and B(36)) xor (A(111) and B(35)) xor (A(112) and B(34)) xor (A(113) and B(33)) xor (A(114) and B(32)) xor (A(115) and B(31)) xor (A(116) and B(30)) xor (A(117) and B(29)) xor (A(118) and B(28)) xor (A(119) and B(27)) xor (A(120) and B(26)) xor (A(121) and B(25)) xor (A(122) and B(24)) xor (A(123) and B(23)) xor (A(124) and B(23)) xor (A(125) and B(21)) xor (A(126) and B(20)) xor (A(20) and B(127)) xor (A(21) and B(126)) xor (A(23) and B(125)) xor (A(23) and B(124)) xor (A(24) and B(123)) xor (A(25) and B(122)) xor (A(26) and B(121)) xor (A(27) and B(120)) xor (A(28) and B(119)) xor (A(29) and B(118)) xor (A(30) and B(117)) xor (A(31) and B(116)) xor (A(32) and B(115)) xor (A(33) and B(114)) xor (A(34) and B(113)) xor (A(35) and B(112)) xor (A(36) and B(111)) xor (A(37) and B(110)) xor (A(38) and B(109)) xor (A(39) and B(108)) xor (A(40) and B(107)) xor (A(41) and B(106)) xor (A(42) and B(105)) xor (A(43) and B(104)) xor (A(44) and B(103)) xor (A(45) and B(102)) xor (A(46) and B(101)) xor (A(47) and B(100)) xor (A(48) and B(99)) xor (A(49) and B(98)) xor (A(50) and B(97)) xor (A(51) and B(96)) xor (A(52) and B(95)) xor (A(53) and B(94)) xor (A(54) and B(93)) xor (A(55) and B(92)) xor (A(56) and B(91)) xor (A(57) and B(90)) xor (A(58) and B(89)) xor (A(59) and B(88)) xor (A(60) and B(87)) xor (A(61) and B(86)) xor (A(62) and B(85)) xor (A(63) and B(84)) xor (A(64) and B(83)) xor (A(65) and B(82)) xor (A(66) and B(81)) xor (A(67) and B(80)) xor (A(68) and B(79)) xor (A(69) and B(78)) xor (A(70) and B(77)) xor (A(71) and B(76)) xor (A(72) and B(75)) xor (A(73) and B(74)) xor (A(74) and B(73)) xor (A(75) and B(72)) xor (A(76) and B(71)) xor (A(77) and B(70)) xor (A(78) and B(69)) xor (A(79) and B(68)) xor (A(80) and B(67)) xor (A(81) and B(66)) xor (A(82) and B(65)) xor (A(83) and B(64)) xor (A(84) and B(63)) xor (A(85) and B(62)) xor (A(86) and B(61)) xor (A(87) and B(60)) xor (A(88) and B(59)) xor (A(89) and B(58)) xor (A(90) and B(57)) xor (A(91) and B(56)) xor (A(92) and B(55)) xor (A(93) and B(54)) xor (A(94) and B(53)) xor (A(95) and B(52)) xor (A(96) and B(51)) xor (A(97) and B(50)) xor (A(98) and B(49)) xor (A(99) and B(48)) xor (A(100) and B(47)) xor (A(101) and B(46)) xor (A(102) and B(45)) xor (A(103) and B(44)) xor (A(104) and B(43)) xor (A(105) and B(42)) xor (A(106) and B(41)) xor (A(107) and B(40)) xor (A(108) and B(39)) xor (A(109) and B(38)) xor (A(110) and B(37)) xor (A(111) and B(36)) xor (A(112) and B(35)) xor (A(113) and B(34)) xor (A(114) and B(33)) xor (A(115) and B(32)) xor (A(116) and B(31)) xor (A(117) and B(30)) xor (A(118) and B(29)) xor (A(119) and B(28)) xor (A(120) and B(27)) xor (A(121) and B(26)) xor (A(122) and B(25)) xor (A(123) and B(24)) xor (A(124) and B(23)) xor (A(125) and B(23)) xor (A(126) and B(22));
    C(21)  <= (A(0) and B(21)) xor (A(1) and B(20)) xor (A(2) and B(19)) xor (A(3) and B(18)) xor (A(4) and B(17)) xor (A(5) and B(16)) xor (A(6) and B(15)) xor (A(7) and B(14)) xor (A(8) and B(13)) xor (A(9) and B(12)) xor (A(10) and B(11)) xor (A(11) and B(10)) xor (A(12) and B(9)) xor (A(13) and B(8)) xor (A(14) and B(7)) xor (A(15) and B(6)) xor (A(16) and B(5)) xor (A(17) and B(4)) xor (A(18) and B(3)) xor (A(19) and B(2)) xor (A(20) and B(1)) xor (A(21) and B(0)) xor (A(14) and B(127)) xor (A(15) and B(126)) xor (A(16) and B(125)) xor (A(17) and B(124)) xor (A(18) and B(123)) xor (A(19) and B(122)) xor (A(20) and B(121)) xor (A(21) and B(120)) xor (A(23) and B(119)) xor (A(23) and B(118)) xor (A(24) and B(117)) xor (A(25) and B(116)) xor (A(26) and B(115)) xor (A(27) and B(114)) xor (A(28) and B(113)) xor (A(29) and B(112)) xor (A(30) and B(111)) xor (A(31) and B(110)) xor (A(32) and B(109)) xor (A(33) and B(108)) xor (A(34) and B(107)) xor (A(35) and B(106)) xor (A(36) and B(105)) xor (A(37) and B(104)) xor (A(38) and B(103)) xor (A(39) and B(102)) xor (A(40) and B(101)) xor (A(41) and B(100)) xor (A(42) and B(99)) xor (A(43) and B(98)) xor (A(44) and B(97)) xor (A(45) and B(96)) xor (A(46) and B(95)) xor (A(47) and B(94)) xor (A(48) and B(93)) xor (A(49) and B(92)) xor (A(50) and B(91)) xor (A(51) and B(90)) xor (A(52) and B(89)) xor (A(53) and B(88)) xor (A(54) and B(87)) xor (A(55) and B(86)) xor (A(56) and B(85)) xor (A(57) and B(84)) xor (A(58) and B(83)) xor (A(59) and B(82)) xor (A(60) and B(81)) xor (A(61) and B(80)) xor (A(62) and B(79)) xor (A(63) and B(78)) xor (A(64) and B(77)) xor (A(65) and B(76)) xor (A(66) and B(75)) xor (A(67) and B(74)) xor (A(68) and B(73)) xor (A(69) and B(72)) xor (A(70) and B(71)) xor (A(71) and B(70)) xor (A(72) and B(69)) xor (A(73) and B(68)) xor (A(74) and B(67)) xor (A(75) and B(66)) xor (A(76) and B(65)) xor (A(77) and B(64)) xor (A(78) and B(63)) xor (A(79) and B(62)) xor (A(80) and B(61)) xor (A(81) and B(60)) xor (A(82) and B(59)) xor (A(83) and B(58)) xor (A(84) and B(57)) xor (A(85) and B(56)) xor (A(86) and B(55)) xor (A(87) and B(54)) xor (A(88) and B(53)) xor (A(89) and B(52)) xor (A(90) and B(51)) xor (A(91) and B(50)) xor (A(92) and B(49)) xor (A(93) and B(48)) xor (A(94) and B(47)) xor (A(95) and B(46)) xor (A(96) and B(45)) xor (A(97) and B(44)) xor (A(98) and B(43)) xor (A(99) and B(42)) xor (A(100) and B(41)) xor (A(101) and B(40)) xor (A(102) and B(39)) xor (A(103) and B(38)) xor (A(104) and B(37)) xor (A(105) and B(36)) xor (A(106) and B(35)) xor (A(107) and B(34)) xor (A(108) and B(33)) xor (A(109) and B(32)) xor (A(110) and B(31)) xor (A(111) and B(30)) xor (A(112) and B(29)) xor (A(113) and B(28)) xor (A(114) and B(27)) xor (A(115) and B(26)) xor (A(116) and B(25)) xor (A(117) and B(24)) xor (A(118) and B(23)) xor (A(119) and B(23)) xor (A(120) and B(21)) xor (A(121) and B(20)) xor (A(122) and B(19)) xor (A(123) and B(18)) xor (A(124) and B(17)) xor (A(125) and B(16)) xor (A(126) and B(15)) xor (A(19) and B(127)) xor (A(20) and B(126)) xor (A(21) and B(125)) xor (A(23) and B(124)) xor (A(23) and B(123)) xor (A(24) and B(122)) xor (A(25) and B(121)) xor (A(26) and B(120)) xor (A(27) and B(119)) xor (A(28) and B(118)) xor (A(29) and B(117)) xor (A(30) and B(116)) xor (A(31) and B(115)) xor (A(32) and B(114)) xor (A(33) and B(113)) xor (A(34) and B(112)) xor (A(35) and B(111)) xor (A(36) and B(110)) xor (A(37) and B(109)) xor (A(38) and B(108)) xor (A(39) and B(107)) xor (A(40) and B(106)) xor (A(41) and B(105)) xor (A(42) and B(104)) xor (A(43) and B(103)) xor (A(44) and B(102)) xor (A(45) and B(101)) xor (A(46) and B(100)) xor (A(47) and B(99)) xor (A(48) and B(98)) xor (A(49) and B(97)) xor (A(50) and B(96)) xor (A(51) and B(95)) xor (A(52) and B(94)) xor (A(53) and B(93)) xor (A(54) and B(92)) xor (A(55) and B(91)) xor (A(56) and B(90)) xor (A(57) and B(89)) xor (A(58) and B(88)) xor (A(59) and B(87)) xor (A(60) and B(86)) xor (A(61) and B(85)) xor (A(62) and B(84)) xor (A(63) and B(83)) xor (A(64) and B(82)) xor (A(65) and B(81)) xor (A(66) and B(80)) xor (A(67) and B(79)) xor (A(68) and B(78)) xor (A(69) and B(77)) xor (A(70) and B(76)) xor (A(71) and B(75)) xor (A(72) and B(74)) xor (A(73) and B(73)) xor (A(74) and B(72)) xor (A(75) and B(71)) xor (A(76) and B(70)) xor (A(77) and B(69)) xor (A(78) and B(68)) xor (A(79) and B(67)) xor (A(80) and B(66)) xor (A(81) and B(65)) xor (A(82) and B(64)) xor (A(83) and B(63)) xor (A(84) and B(62)) xor (A(85) and B(61)) xor (A(86) and B(60)) xor (A(87) and B(59)) xor (A(88) and B(58)) xor (A(89) and B(57)) xor (A(90) and B(56)) xor (A(91) and B(55)) xor (A(92) and B(54)) xor (A(93) and B(53)) xor (A(94) and B(52)) xor (A(95) and B(51)) xor (A(96) and B(50)) xor (A(97) and B(49)) xor (A(98) and B(48)) xor (A(99) and B(47)) xor (A(100) and B(46)) xor (A(101) and B(45)) xor (A(102) and B(44)) xor (A(103) and B(43)) xor (A(104) and B(42)) xor (A(105) and B(41)) xor (A(106) and B(40)) xor (A(107) and B(39)) xor (A(108) and B(38)) xor (A(109) and B(37)) xor (A(110) and B(36)) xor (A(111) and B(35)) xor (A(112) and B(34)) xor (A(113) and B(33)) xor (A(114) and B(32)) xor (A(115) and B(31)) xor (A(116) and B(30)) xor (A(117) and B(29)) xor (A(118) and B(28)) xor (A(119) and B(27)) xor (A(120) and B(26)) xor (A(121) and B(25)) xor (A(122) and B(24)) xor (A(123) and B(23)) xor (A(124) and B(23)) xor (A(125) and B(21)) xor (A(126) and B(20)) xor (A(20) and B(127)) xor (A(21) and B(126)) xor (A(23) and B(125)) xor (A(23) and B(124)) xor (A(24) and B(123)) xor (A(25) and B(122)) xor (A(26) and B(121)) xor (A(27) and B(120)) xor (A(28) and B(119)) xor (A(29) and B(118)) xor (A(30) and B(117)) xor (A(31) and B(116)) xor (A(32) and B(115)) xor (A(33) and B(114)) xor (A(34) and B(113)) xor (A(35) and B(112)) xor (A(36) and B(111)) xor (A(37) and B(110)) xor (A(38) and B(109)) xor (A(39) and B(108)) xor (A(40) and B(107)) xor (A(41) and B(106)) xor (A(42) and B(105)) xor (A(43) and B(104)) xor (A(44) and B(103)) xor (A(45) and B(102)) xor (A(46) and B(101)) xor (A(47) and B(100)) xor (A(48) and B(99)) xor (A(49) and B(98)) xor (A(50) and B(97)) xor (A(51) and B(96)) xor (A(52) and B(95)) xor (A(53) and B(94)) xor (A(54) and B(93)) xor (A(55) and B(92)) xor (A(56) and B(91)) xor (A(57) and B(90)) xor (A(58) and B(89)) xor (A(59) and B(88)) xor (A(60) and B(87)) xor (A(61) and B(86)) xor (A(62) and B(85)) xor (A(63) and B(84)) xor (A(64) and B(83)) xor (A(65) and B(82)) xor (A(66) and B(81)) xor (A(67) and B(80)) xor (A(68) and B(79)) xor (A(69) and B(78)) xor (A(70) and B(77)) xor (A(71) and B(76)) xor (A(72) and B(75)) xor (A(73) and B(74)) xor (A(74) and B(73)) xor (A(75) and B(72)) xor (A(76) and B(71)) xor (A(77) and B(70)) xor (A(78) and B(69)) xor (A(79) and B(68)) xor (A(80) and B(67)) xor (A(81) and B(66)) xor (A(82) and B(65)) xor (A(83) and B(64)) xor (A(84) and B(63)) xor (A(85) and B(62)) xor (A(86) and B(61)) xor (A(87) and B(60)) xor (A(88) and B(59)) xor (A(89) and B(58)) xor (A(90) and B(57)) xor (A(91) and B(56)) xor (A(92) and B(55)) xor (A(93) and B(54)) xor (A(94) and B(53)) xor (A(95) and B(52)) xor (A(96) and B(51)) xor (A(97) and B(50)) xor (A(98) and B(49)) xor (A(99) and B(48)) xor (A(100) and B(47)) xor (A(101) and B(46)) xor (A(102) and B(45)) xor (A(103) and B(44)) xor (A(104) and B(43)) xor (A(105) and B(42)) xor (A(106) and B(41)) xor (A(107) and B(40)) xor (A(108) and B(39)) xor (A(109) and B(38)) xor (A(110) and B(37)) xor (A(111) and B(36)) xor (A(112) and B(35)) xor (A(113) and B(34)) xor (A(114) and B(33)) xor (A(115) and B(32)) xor (A(116) and B(31)) xor (A(117) and B(30)) xor (A(118) and B(29)) xor (A(119) and B(28)) xor (A(120) and B(27)) xor (A(121) and B(26)) xor (A(122) and B(25)) xor (A(123) and B(24)) xor (A(124) and B(23)) xor (A(125) and B(23)) xor (A(126) and B(21)) xor (A(21) and B(127)) xor (A(23) and B(126)) xor (A(23) and B(125)) xor (A(24) and B(124)) xor (A(25) and B(123)) xor (A(26) and B(122)) xor (A(27) and B(121)) xor (A(28) and B(120)) xor (A(29) and B(119)) xor (A(30) and B(118)) xor (A(31) and B(117)) xor (A(32) and B(116)) xor (A(33) and B(115)) xor (A(34) and B(114)) xor (A(35) and B(113)) xor (A(36) and B(112)) xor (A(37) and B(111)) xor (A(38) and B(110)) xor (A(39) and B(109)) xor (A(40) and B(108)) xor (A(41) and B(107)) xor (A(42) and B(106)) xor (A(43) and B(105)) xor (A(44) and B(104)) xor (A(45) and B(103)) xor (A(46) and B(102)) xor (A(47) and B(101)) xor (A(48) and B(100)) xor (A(49) and B(99)) xor (A(50) and B(98)) xor (A(51) and B(97)) xor (A(52) and B(96)) xor (A(53) and B(95)) xor (A(54) and B(94)) xor (A(55) and B(93)) xor (A(56) and B(92)) xor (A(57) and B(91)) xor (A(58) and B(90)) xor (A(59) and B(89)) xor (A(60) and B(88)) xor (A(61) and B(87)) xor (A(62) and B(86)) xor (A(63) and B(85)) xor (A(64) and B(84)) xor (A(65) and B(83)) xor (A(66) and B(82)) xor (A(67) and B(81)) xor (A(68) and B(80)) xor (A(69) and B(79)) xor (A(70) and B(78)) xor (A(71) and B(77)) xor (A(72) and B(76)) xor (A(73) and B(75)) xor (A(74) and B(74)) xor (A(75) and B(73)) xor (A(76) and B(72)) xor (A(77) and B(71)) xor (A(78) and B(70)) xor (A(79) and B(69)) xor (A(80) and B(68)) xor (A(81) and B(67)) xor (A(82) and B(66)) xor (A(83) and B(65)) xor (A(84) and B(64)) xor (A(85) and B(63)) xor (A(86) and B(62)) xor (A(87) and B(61)) xor (A(88) and B(60)) xor (A(89) and B(59)) xor (A(90) and B(58)) xor (A(91) and B(57)) xor (A(92) and B(56)) xor (A(93) and B(55)) xor (A(94) and B(54)) xor (A(95) and B(53)) xor (A(96) and B(52)) xor (A(97) and B(51)) xor (A(98) and B(50)) xor (A(99) and B(49)) xor (A(100) and B(48)) xor (A(101) and B(47)) xor (A(102) and B(46)) xor (A(103) and B(45)) xor (A(104) and B(44)) xor (A(105) and B(43)) xor (A(106) and B(42)) xor (A(107) and B(41)) xor (A(108) and B(40)) xor (A(109) and B(39)) xor (A(110) and B(38)) xor (A(111) and B(37)) xor (A(112) and B(36)) xor (A(113) and B(35)) xor (A(114) and B(34)) xor (A(115) and B(33)) xor (A(116) and B(32)) xor (A(117) and B(31)) xor (A(118) and B(30)) xor (A(119) and B(29)) xor (A(120) and B(28)) xor (A(121) and B(27)) xor (A(122) and B(26)) xor (A(123) and B(25)) xor (A(124) and B(24)) xor (A(125) and B(23)) xor (A(126) and B(23));
    C(22)  <= (A(0) and B(23)) xor (A(1) and B(21)) xor (A(2) and B(20)) xor (A(3) and B(19)) xor (A(4) and B(18)) xor (A(5) and B(17)) xor (A(6) and B(16)) xor (A(7) and B(15)) xor (A(8) and B(14)) xor (A(9) and B(13)) xor (A(10) and B(12)) xor (A(11) and B(11)) xor (A(12) and B(10)) xor (A(13) and B(9)) xor (A(14) and B(8)) xor (A(15) and B(7)) xor (A(16) and B(6)) xor (A(17) and B(5)) xor (A(18) and B(4)) xor (A(19) and B(3)) xor (A(20) and B(2)) xor (A(21) and B(1)) xor (A(23) and B(0)) xor (A(15) and B(127)) xor (A(16) and B(126)) xor (A(17) and B(125)) xor (A(18) and B(124)) xor (A(19) and B(123)) xor (A(20) and B(122)) xor (A(21) and B(121)) xor (A(23) and B(120)) xor (A(23) and B(119)) xor (A(24) and B(118)) xor (A(25) and B(117)) xor (A(26) and B(116)) xor (A(27) and B(115)) xor (A(28) and B(114)) xor (A(29) and B(113)) xor (A(30) and B(112)) xor (A(31) and B(111)) xor (A(32) and B(110)) xor (A(33) and B(109)) xor (A(34) and B(108)) xor (A(35) and B(107)) xor (A(36) and B(106)) xor (A(37) and B(105)) xor (A(38) and B(104)) xor (A(39) and B(103)) xor (A(40) and B(102)) xor (A(41) and B(101)) xor (A(42) and B(100)) xor (A(43) and B(99)) xor (A(44) and B(98)) xor (A(45) and B(97)) xor (A(46) and B(96)) xor (A(47) and B(95)) xor (A(48) and B(94)) xor (A(49) and B(93)) xor (A(50) and B(92)) xor (A(51) and B(91)) xor (A(52) and B(90)) xor (A(53) and B(89)) xor (A(54) and B(88)) xor (A(55) and B(87)) xor (A(56) and B(86)) xor (A(57) and B(85)) xor (A(58) and B(84)) xor (A(59) and B(83)) xor (A(60) and B(82)) xor (A(61) and B(81)) xor (A(62) and B(80)) xor (A(63) and B(79)) xor (A(64) and B(78)) xor (A(65) and B(77)) xor (A(66) and B(76)) xor (A(67) and B(75)) xor (A(68) and B(74)) xor (A(69) and B(73)) xor (A(70) and B(72)) xor (A(71) and B(71)) xor (A(72) and B(70)) xor (A(73) and B(69)) xor (A(74) and B(68)) xor (A(75) and B(67)) xor (A(76) and B(66)) xor (A(77) and B(65)) xor (A(78) and B(64)) xor (A(79) and B(63)) xor (A(80) and B(62)) xor (A(81) and B(61)) xor (A(82) and B(60)) xor (A(83) and B(59)) xor (A(84) and B(58)) xor (A(85) and B(57)) xor (A(86) and B(56)) xor (A(87) and B(55)) xor (A(88) and B(54)) xor (A(89) and B(53)) xor (A(90) and B(52)) xor (A(91) and B(51)) xor (A(92) and B(50)) xor (A(93) and B(49)) xor (A(94) and B(48)) xor (A(95) and B(47)) xor (A(96) and B(46)) xor (A(97) and B(45)) xor (A(98) and B(44)) xor (A(99) and B(43)) xor (A(100) and B(42)) xor (A(101) and B(41)) xor (A(102) and B(40)) xor (A(103) and B(39)) xor (A(104) and B(38)) xor (A(105) and B(37)) xor (A(106) and B(36)) xor (A(107) and B(35)) xor (A(108) and B(34)) xor (A(109) and B(33)) xor (A(110) and B(32)) xor (A(111) and B(31)) xor (A(112) and B(30)) xor (A(113) and B(29)) xor (A(114) and B(28)) xor (A(115) and B(27)) xor (A(116) and B(26)) xor (A(117) and B(25)) xor (A(118) and B(24)) xor (A(119) and B(23)) xor (A(120) and B(23)) xor (A(121) and B(21)) xor (A(122) and B(20)) xor (A(123) and B(19)) xor (A(124) and B(18)) xor (A(125) and B(17)) xor (A(126) and B(16)) xor (A(20) and B(127)) xor (A(21) and B(126)) xor (A(23) and B(125)) xor (A(23) and B(124)) xor (A(24) and B(123)) xor (A(25) and B(122)) xor (A(26) and B(121)) xor (A(27) and B(120)) xor (A(28) and B(119)) xor (A(29) and B(118)) xor (A(30) and B(117)) xor (A(31) and B(116)) xor (A(32) and B(115)) xor (A(33) and B(114)) xor (A(34) and B(113)) xor (A(35) and B(112)) xor (A(36) and B(111)) xor (A(37) and B(110)) xor (A(38) and B(109)) xor (A(39) and B(108)) xor (A(40) and B(107)) xor (A(41) and B(106)) xor (A(42) and B(105)) xor (A(43) and B(104)) xor (A(44) and B(103)) xor (A(45) and B(102)) xor (A(46) and B(101)) xor (A(47) and B(100)) xor (A(48) and B(99)) xor (A(49) and B(98)) xor (A(50) and B(97)) xor (A(51) and B(96)) xor (A(52) and B(95)) xor (A(53) and B(94)) xor (A(54) and B(93)) xor (A(55) and B(92)) xor (A(56) and B(91)) xor (A(57) and B(90)) xor (A(58) and B(89)) xor (A(59) and B(88)) xor (A(60) and B(87)) xor (A(61) and B(86)) xor (A(62) and B(85)) xor (A(63) and B(84)) xor (A(64) and B(83)) xor (A(65) and B(82)) xor (A(66) and B(81)) xor (A(67) and B(80)) xor (A(68) and B(79)) xor (A(69) and B(78)) xor (A(70) and B(77)) xor (A(71) and B(76)) xor (A(72) and B(75)) xor (A(73) and B(74)) xor (A(74) and B(73)) xor (A(75) and B(72)) xor (A(76) and B(71)) xor (A(77) and B(70)) xor (A(78) and B(69)) xor (A(79) and B(68)) xor (A(80) and B(67)) xor (A(81) and B(66)) xor (A(82) and B(65)) xor (A(83) and B(64)) xor (A(84) and B(63)) xor (A(85) and B(62)) xor (A(86) and B(61)) xor (A(87) and B(60)) xor (A(88) and B(59)) xor (A(89) and B(58)) xor (A(90) and B(57)) xor (A(91) and B(56)) xor (A(92) and B(55)) xor (A(93) and B(54)) xor (A(94) and B(53)) xor (A(95) and B(52)) xor (A(96) and B(51)) xor (A(97) and B(50)) xor (A(98) and B(49)) xor (A(99) and B(48)) xor (A(100) and B(47)) xor (A(101) and B(46)) xor (A(102) and B(45)) xor (A(103) and B(44)) xor (A(104) and B(43)) xor (A(105) and B(42)) xor (A(106) and B(41)) xor (A(107) and B(40)) xor (A(108) and B(39)) xor (A(109) and B(38)) xor (A(110) and B(37)) xor (A(111) and B(36)) xor (A(112) and B(35)) xor (A(113) and B(34)) xor (A(114) and B(33)) xor (A(115) and B(32)) xor (A(116) and B(31)) xor (A(117) and B(30)) xor (A(118) and B(29)) xor (A(119) and B(28)) xor (A(120) and B(27)) xor (A(121) and B(26)) xor (A(122) and B(25)) xor (A(123) and B(24)) xor (A(124) and B(23)) xor (A(125) and B(23)) xor (A(126) and B(21)) xor (A(21) and B(127)) xor (A(23) and B(126)) xor (A(23) and B(125)) xor (A(24) and B(124)) xor (A(25) and B(123)) xor (A(26) and B(122)) xor (A(27) and B(121)) xor (A(28) and B(120)) xor (A(29) and B(119)) xor (A(30) and B(118)) xor (A(31) and B(117)) xor (A(32) and B(116)) xor (A(33) and B(115)) xor (A(34) and B(114)) xor (A(35) and B(113)) xor (A(36) and B(112)) xor (A(37) and B(111)) xor (A(38) and B(110)) xor (A(39) and B(109)) xor (A(40) and B(108)) xor (A(41) and B(107)) xor (A(42) and B(106)) xor (A(43) and B(105)) xor (A(44) and B(104)) xor (A(45) and B(103)) xor (A(46) and B(102)) xor (A(47) and B(101)) xor (A(48) and B(100)) xor (A(49) and B(99)) xor (A(50) and B(98)) xor (A(51) and B(97)) xor (A(52) and B(96)) xor (A(53) and B(95)) xor (A(54) and B(94)) xor (A(55) and B(93)) xor (A(56) and B(92)) xor (A(57) and B(91)) xor (A(58) and B(90)) xor (A(59) and B(89)) xor (A(60) and B(88)) xor (A(61) and B(87)) xor (A(62) and B(86)) xor (A(63) and B(85)) xor (A(64) and B(84)) xor (A(65) and B(83)) xor (A(66) and B(82)) xor (A(67) and B(81)) xor (A(68) and B(80)) xor (A(69) and B(79)) xor (A(70) and B(78)) xor (A(71) and B(77)) xor (A(72) and B(76)) xor (A(73) and B(75)) xor (A(74) and B(74)) xor (A(75) and B(73)) xor (A(76) and B(72)) xor (A(77) and B(71)) xor (A(78) and B(70)) xor (A(79) and B(69)) xor (A(80) and B(68)) xor (A(81) and B(67)) xor (A(82) and B(66)) xor (A(83) and B(65)) xor (A(84) and B(64)) xor (A(85) and B(63)) xor (A(86) and B(62)) xor (A(87) and B(61)) xor (A(88) and B(60)) xor (A(89) and B(59)) xor (A(90) and B(58)) xor (A(91) and B(57)) xor (A(92) and B(56)) xor (A(93) and B(55)) xor (A(94) and B(54)) xor (A(95) and B(53)) xor (A(96) and B(52)) xor (A(97) and B(51)) xor (A(98) and B(50)) xor (A(99) and B(49)) xor (A(100) and B(48)) xor (A(101) and B(47)) xor (A(102) and B(46)) xor (A(103) and B(45)) xor (A(104) and B(44)) xor (A(105) and B(43)) xor (A(106) and B(42)) xor (A(107) and B(41)) xor (A(108) and B(40)) xor (A(109) and B(39)) xor (A(110) and B(38)) xor (A(111) and B(37)) xor (A(112) and B(36)) xor (A(113) and B(35)) xor (A(114) and B(34)) xor (A(115) and B(33)) xor (A(116) and B(32)) xor (A(117) and B(31)) xor (A(118) and B(30)) xor (A(119) and B(29)) xor (A(120) and B(28)) xor (A(121) and B(27)) xor (A(122) and B(26)) xor (A(123) and B(25)) xor (A(124) and B(24)) xor (A(125) and B(23)) xor (A(126) and B(23)) xor (A(23) and B(127)) xor (A(23) and B(126)) xor (A(24) and B(125)) xor (A(25) and B(124)) xor (A(26) and B(123)) xor (A(27) and B(122)) xor (A(28) and B(121)) xor (A(29) and B(120)) xor (A(30) and B(119)) xor (A(31) and B(118)) xor (A(32) and B(117)) xor (A(33) and B(116)) xor (A(34) and B(115)) xor (A(35) and B(114)) xor (A(36) and B(113)) xor (A(37) and B(112)) xor (A(38) and B(111)) xor (A(39) and B(110)) xor (A(40) and B(109)) xor (A(41) and B(108)) xor (A(42) and B(107)) xor (A(43) and B(106)) xor (A(44) and B(105)) xor (A(45) and B(104)) xor (A(46) and B(103)) xor (A(47) and B(102)) xor (A(48) and B(101)) xor (A(49) and B(100)) xor (A(50) and B(99)) xor (A(51) and B(98)) xor (A(52) and B(97)) xor (A(53) and B(96)) xor (A(54) and B(95)) xor (A(55) and B(94)) xor (A(56) and B(93)) xor (A(57) and B(92)) xor (A(58) and B(91)) xor (A(59) and B(90)) xor (A(60) and B(89)) xor (A(61) and B(88)) xor (A(62) and B(87)) xor (A(63) and B(86)) xor (A(64) and B(85)) xor (A(65) and B(84)) xor (A(66) and B(83)) xor (A(67) and B(82)) xor (A(68) and B(81)) xor (A(69) and B(80)) xor (A(70) and B(79)) xor (A(71) and B(78)) xor (A(72) and B(77)) xor (A(73) and B(76)) xor (A(74) and B(75)) xor (A(75) and B(74)) xor (A(76) and B(73)) xor (A(77) and B(72)) xor (A(78) and B(71)) xor (A(79) and B(70)) xor (A(80) and B(69)) xor (A(81) and B(68)) xor (A(82) and B(67)) xor (A(83) and B(66)) xor (A(84) and B(65)) xor (A(85) and B(64)) xor (A(86) and B(63)) xor (A(87) and B(62)) xor (A(88) and B(61)) xor (A(89) and B(60)) xor (A(90) and B(59)) xor (A(91) and B(58)) xor (A(92) and B(57)) xor (A(93) and B(56)) xor (A(94) and B(55)) xor (A(95) and B(54)) xor (A(96) and B(53)) xor (A(97) and B(52)) xor (A(98) and B(51)) xor (A(99) and B(50)) xor (A(100) and B(49)) xor (A(101) and B(48)) xor (A(102) and B(47)) xor (A(103) and B(46)) xor (A(104) and B(45)) xor (A(105) and B(44)) xor (A(106) and B(43)) xor (A(107) and B(42)) xor (A(108) and B(41)) xor (A(109) and B(40)) xor (A(110) and B(39)) xor (A(111) and B(38)) xor (A(112) and B(37)) xor (A(113) and B(36)) xor (A(114) and B(35)) xor (A(115) and B(34)) xor (A(116) and B(33)) xor (A(117) and B(32)) xor (A(118) and B(31)) xor (A(119) and B(30)) xor (A(120) and B(29)) xor (A(121) and B(28)) xor (A(122) and B(27)) xor (A(123) and B(26)) xor (A(124) and B(25)) xor (A(125) and B(24)) xor (A(126) and B(24));
    C(23)  <= (A(0) and B(23)) xor (A(1) and B(23)) xor (A(2) and B(21)) xor (A(3) and B(20)) xor (A(4) and B(19)) xor (A(5) and B(18)) xor (A(6) and B(17)) xor (A(7) and B(16)) xor (A(8) and B(15)) xor (A(9) and B(14)) xor (A(10) and B(13)) xor (A(11) and B(12)) xor (A(12) and B(11)) xor (A(13) and B(10)) xor (A(14) and B(9)) xor (A(15) and B(8)) xor (A(16) and B(7)) xor (A(17) and B(6)) xor (A(18) and B(5)) xor (A(19) and B(4)) xor (A(20) and B(3)) xor (A(21) and B(2)) xor (A(23) and B(1)) xor (A(23) and B(0)) xor (A(16) and B(127)) xor (A(17) and B(126)) xor (A(18) and B(125)) xor (A(19) and B(124)) xor (A(20) and B(123)) xor (A(21) and B(122)) xor (A(23) and B(121)) xor (A(23) and B(120)) xor (A(24) and B(119)) xor (A(25) and B(118)) xor (A(26) and B(117)) xor (A(27) and B(116)) xor (A(28) and B(115)) xor (A(29) and B(114)) xor (A(30) and B(113)) xor (A(31) and B(112)) xor (A(32) and B(111)) xor (A(33) and B(110)) xor (A(34) and B(109)) xor (A(35) and B(108)) xor (A(36) and B(107)) xor (A(37) and B(106)) xor (A(38) and B(105)) xor (A(39) and B(104)) xor (A(40) and B(103)) xor (A(41) and B(102)) xor (A(42) and B(101)) xor (A(43) and B(100)) xor (A(44) and B(99)) xor (A(45) and B(98)) xor (A(46) and B(97)) xor (A(47) and B(96)) xor (A(48) and B(95)) xor (A(49) and B(94)) xor (A(50) and B(93)) xor (A(51) and B(92)) xor (A(52) and B(91)) xor (A(53) and B(90)) xor (A(54) and B(89)) xor (A(55) and B(88)) xor (A(56) and B(87)) xor (A(57) and B(86)) xor (A(58) and B(85)) xor (A(59) and B(84)) xor (A(60) and B(83)) xor (A(61) and B(82)) xor (A(62) and B(81)) xor (A(63) and B(80)) xor (A(64) and B(79)) xor (A(65) and B(78)) xor (A(66) and B(77)) xor (A(67) and B(76)) xor (A(68) and B(75)) xor (A(69) and B(74)) xor (A(70) and B(73)) xor (A(71) and B(72)) xor (A(72) and B(71)) xor (A(73) and B(70)) xor (A(74) and B(69)) xor (A(75) and B(68)) xor (A(76) and B(67)) xor (A(77) and B(66)) xor (A(78) and B(65)) xor (A(79) and B(64)) xor (A(80) and B(63)) xor (A(81) and B(62)) xor (A(82) and B(61)) xor (A(83) and B(60)) xor (A(84) and B(59)) xor (A(85) and B(58)) xor (A(86) and B(57)) xor (A(87) and B(56)) xor (A(88) and B(55)) xor (A(89) and B(54)) xor (A(90) and B(53)) xor (A(91) and B(52)) xor (A(92) and B(51)) xor (A(93) and B(50)) xor (A(94) and B(49)) xor (A(95) and B(48)) xor (A(96) and B(47)) xor (A(97) and B(46)) xor (A(98) and B(45)) xor (A(99) and B(44)) xor (A(100) and B(43)) xor (A(101) and B(42)) xor (A(102) and B(41)) xor (A(103) and B(40)) xor (A(104) and B(39)) xor (A(105) and B(38)) xor (A(106) and B(37)) xor (A(107) and B(36)) xor (A(108) and B(35)) xor (A(109) and B(34)) xor (A(110) and B(33)) xor (A(111) and B(32)) xor (A(112) and B(31)) xor (A(113) and B(30)) xor (A(114) and B(29)) xor (A(115) and B(28)) xor (A(116) and B(27)) xor (A(117) and B(26)) xor (A(118) and B(25)) xor (A(119) and B(24)) xor (A(120) and B(23)) xor (A(121) and B(23)) xor (A(122) and B(21)) xor (A(123) and B(20)) xor (A(124) and B(19)) xor (A(125) and B(18)) xor (A(126) and B(17)) xor (A(21) and B(127)) xor (A(23) and B(126)) xor (A(23) and B(125)) xor (A(24) and B(124)) xor (A(25) and B(123)) xor (A(26) and B(122)) xor (A(27) and B(121)) xor (A(28) and B(120)) xor (A(29) and B(119)) xor (A(30) and B(118)) xor (A(31) and B(117)) xor (A(32) and B(116)) xor (A(33) and B(115)) xor (A(34) and B(114)) xor (A(35) and B(113)) xor (A(36) and B(112)) xor (A(37) and B(111)) xor (A(38) and B(110)) xor (A(39) and B(109)) xor (A(40) and B(108)) xor (A(41) and B(107)) xor (A(42) and B(106)) xor (A(43) and B(105)) xor (A(44) and B(104)) xor (A(45) and B(103)) xor (A(46) and B(102)) xor (A(47) and B(101)) xor (A(48) and B(100)) xor (A(49) and B(99)) xor (A(50) and B(98)) xor (A(51) and B(97)) xor (A(52) and B(96)) xor (A(53) and B(95)) xor (A(54) and B(94)) xor (A(55) and B(93)) xor (A(56) and B(92)) xor (A(57) and B(91)) xor (A(58) and B(90)) xor (A(59) and B(89)) xor (A(60) and B(88)) xor (A(61) and B(87)) xor (A(62) and B(86)) xor (A(63) and B(85)) xor (A(64) and B(84)) xor (A(65) and B(83)) xor (A(66) and B(82)) xor (A(67) and B(81)) xor (A(68) and B(80)) xor (A(69) and B(79)) xor (A(70) and B(78)) xor (A(71) and B(77)) xor (A(72) and B(76)) xor (A(73) and B(75)) xor (A(74) and B(74)) xor (A(75) and B(73)) xor (A(76) and B(72)) xor (A(77) and B(71)) xor (A(78) and B(70)) xor (A(79) and B(69)) xor (A(80) and B(68)) xor (A(81) and B(67)) xor (A(82) and B(66)) xor (A(83) and B(65)) xor (A(84) and B(64)) xor (A(85) and B(63)) xor (A(86) and B(62)) xor (A(87) and B(61)) xor (A(88) and B(60)) xor (A(89) and B(59)) xor (A(90) and B(58)) xor (A(91) and B(57)) xor (A(92) and B(56)) xor (A(93) and B(55)) xor (A(94) and B(54)) xor (A(95) and B(53)) xor (A(96) and B(52)) xor (A(97) and B(51)) xor (A(98) and B(50)) xor (A(99) and B(49)) xor (A(100) and B(48)) xor (A(101) and B(47)) xor (A(102) and B(46)) xor (A(103) and B(45)) xor (A(104) and B(44)) xor (A(105) and B(43)) xor (A(106) and B(42)) xor (A(107) and B(41)) xor (A(108) and B(40)) xor (A(109) and B(39)) xor (A(110) and B(38)) xor (A(111) and B(37)) xor (A(112) and B(36)) xor (A(113) and B(35)) xor (A(114) and B(34)) xor (A(115) and B(33)) xor (A(116) and B(32)) xor (A(117) and B(31)) xor (A(118) and B(30)) xor (A(119) and B(29)) xor (A(120) and B(28)) xor (A(121) and B(27)) xor (A(122) and B(26)) xor (A(123) and B(25)) xor (A(124) and B(24)) xor (A(125) and B(23)) xor (A(126) and B(23)) xor (A(23) and B(127)) xor (A(23) and B(126)) xor (A(24) and B(125)) xor (A(25) and B(124)) xor (A(26) and B(123)) xor (A(27) and B(122)) xor (A(28) and B(121)) xor (A(29) and B(120)) xor (A(30) and B(119)) xor (A(31) and B(118)) xor (A(32) and B(117)) xor (A(33) and B(116)) xor (A(34) and B(115)) xor (A(35) and B(114)) xor (A(36) and B(113)) xor (A(37) and B(112)) xor (A(38) and B(111)) xor (A(39) and B(110)) xor (A(40) and B(109)) xor (A(41) and B(108)) xor (A(42) and B(107)) xor (A(43) and B(106)) xor (A(44) and B(105)) xor (A(45) and B(104)) xor (A(46) and B(103)) xor (A(47) and B(102)) xor (A(48) and B(101)) xor (A(49) and B(100)) xor (A(50) and B(99)) xor (A(51) and B(98)) xor (A(52) and B(97)) xor (A(53) and B(96)) xor (A(54) and B(95)) xor (A(55) and B(94)) xor (A(56) and B(93)) xor (A(57) and B(92)) xor (A(58) and B(91)) xor (A(59) and B(90)) xor (A(60) and B(89)) xor (A(61) and B(88)) xor (A(62) and B(87)) xor (A(63) and B(86)) xor (A(64) and B(85)) xor (A(65) and B(84)) xor (A(66) and B(83)) xor (A(67) and B(82)) xor (A(68) and B(81)) xor (A(69) and B(80)) xor (A(70) and B(79)) xor (A(71) and B(78)) xor (A(72) and B(77)) xor (A(73) and B(76)) xor (A(74) and B(75)) xor (A(75) and B(74)) xor (A(76) and B(73)) xor (A(77) and B(72)) xor (A(78) and B(71)) xor (A(79) and B(70)) xor (A(80) and B(69)) xor (A(81) and B(68)) xor (A(82) and B(67)) xor (A(83) and B(66)) xor (A(84) and B(65)) xor (A(85) and B(64)) xor (A(86) and B(63)) xor (A(87) and B(62)) xor (A(88) and B(61)) xor (A(89) and B(60)) xor (A(90) and B(59)) xor (A(91) and B(58)) xor (A(92) and B(57)) xor (A(93) and B(56)) xor (A(94) and B(55)) xor (A(95) and B(54)) xor (A(96) and B(53)) xor (A(97) and B(52)) xor (A(98) and B(51)) xor (A(99) and B(50)) xor (A(100) and B(49)) xor (A(101) and B(48)) xor (A(102) and B(47)) xor (A(103) and B(46)) xor (A(104) and B(45)) xor (A(105) and B(44)) xor (A(106) and B(43)) xor (A(107) and B(42)) xor (A(108) and B(41)) xor (A(109) and B(40)) xor (A(110) and B(39)) xor (A(111) and B(38)) xor (A(112) and B(37)) xor (A(113) and B(36)) xor (A(114) and B(35)) xor (A(115) and B(34)) xor (A(116) and B(33)) xor (A(117) and B(32)) xor (A(118) and B(31)) xor (A(119) and B(30)) xor (A(120) and B(29)) xor (A(121) and B(28)) xor (A(122) and B(27)) xor (A(123) and B(26)) xor (A(124) and B(25)) xor (A(125) and B(24)) xor (A(126) and B(23)) xor (A(23) and B(127)) xor (A(24) and B(126)) xor (A(25) and B(125)) xor (A(26) and B(124)) xor (A(27) and B(123)) xor (A(28) and B(122)) xor (A(29) and B(121)) xor (A(30) and B(120)) xor (A(31) and B(119)) xor (A(32) and B(118)) xor (A(33) and B(117)) xor (A(34) and B(116)) xor (A(35) and B(115)) xor (A(36) and B(114)) xor (A(37) and B(113)) xor (A(38) and B(112)) xor (A(39) and B(111)) xor (A(40) and B(110)) xor (A(41) and B(109)) xor (A(42) and B(108)) xor (A(43) and B(107)) xor (A(44) and B(106)) xor (A(45) and B(105)) xor (A(46) and B(104)) xor (A(47) and B(103)) xor (A(48) and B(102)) xor (A(49) and B(101)) xor (A(50) and B(100)) xor (A(51) and B(99)) xor (A(52) and B(98)) xor (A(53) and B(97)) xor (A(54) and B(96)) xor (A(55) and B(95)) xor (A(56) and B(94)) xor (A(57) and B(93)) xor (A(58) and B(92)) xor (A(59) and B(91)) xor (A(60) and B(90)) xor (A(61) and B(89)) xor (A(62) and B(88)) xor (A(63) and B(87)) xor (A(64) and B(86)) xor (A(65) and B(85)) xor (A(66) and B(84)) xor (A(67) and B(83)) xor (A(68) and B(82)) xor (A(69) and B(81)) xor (A(70) and B(80)) xor (A(71) and B(79)) xor (A(72) and B(78)) xor (A(73) and B(77)) xor (A(74) and B(76)) xor (A(75) and B(75)) xor (A(76) and B(74)) xor (A(77) and B(73)) xor (A(78) and B(72)) xor (A(79) and B(71)) xor (A(80) and B(70)) xor (A(81) and B(69)) xor (A(82) and B(68)) xor (A(83) and B(67)) xor (A(84) and B(66)) xor (A(85) and B(65)) xor (A(86) and B(64)) xor (A(87) and B(63)) xor (A(88) and B(62)) xor (A(89) and B(61)) xor (A(90) and B(60)) xor (A(91) and B(59)) xor (A(92) and B(58)) xor (A(93) and B(57)) xor (A(94) and B(56)) xor (A(95) and B(55)) xor (A(96) and B(54)) xor (A(97) and B(53)) xor (A(98) and B(52)) xor (A(99) and B(51)) xor (A(100) and B(50)) xor (A(101) and B(49)) xor (A(102) and B(48)) xor (A(103) and B(47)) xor (A(104) and B(46)) xor (A(105) and B(45)) xor (A(106) and B(44)) xor (A(107) and B(43)) xor (A(108) and B(42)) xor (A(109) and B(41)) xor (A(110) and B(40)) xor (A(111) and B(39)) xor (A(112) and B(38)) xor (A(113) and B(37)) xor (A(114) and B(36)) xor (A(115) and B(35)) xor (A(116) and B(34)) xor (A(117) and B(33)) xor (A(118) and B(32)) xor (A(119) and B(31)) xor (A(120) and B(30)) xor (A(121) and B(29)) xor (A(122) and B(28)) xor (A(123) and B(27)) xor (A(124) and B(26)) xor (A(125) and B(25)) xor (A(126) and B(25));
    C(24)  <= (A(0) and B(24)) xor (A(1) and B(23)) xor (A(2) and B(23)) xor (A(3) and B(21)) xor (A(4) and B(20)) xor (A(5) and B(19)) xor (A(6) and B(18)) xor (A(7) and B(17)) xor (A(8) and B(16)) xor (A(9) and B(15)) xor (A(10) and B(14)) xor (A(11) and B(13)) xor (A(12) and B(12)) xor (A(13) and B(11)) xor (A(14) and B(10)) xor (A(15) and B(9)) xor (A(16) and B(8)) xor (A(17) and B(7)) xor (A(18) and B(6)) xor (A(19) and B(5)) xor (A(20) and B(4)) xor (A(21) and B(3)) xor (A(23) and B(2)) xor (A(23) and B(1)) xor (A(24) and B(0)) xor (A(17) and B(127)) xor (A(18) and B(126)) xor (A(19) and B(125)) xor (A(20) and B(124)) xor (A(21) and B(123)) xor (A(23) and B(122)) xor (A(23) and B(121)) xor (A(24) and B(120)) xor (A(25) and B(119)) xor (A(26) and B(118)) xor (A(27) and B(117)) xor (A(28) and B(116)) xor (A(29) and B(115)) xor (A(30) and B(114)) xor (A(31) and B(113)) xor (A(32) and B(112)) xor (A(33) and B(111)) xor (A(34) and B(110)) xor (A(35) and B(109)) xor (A(36) and B(108)) xor (A(37) and B(107)) xor (A(38) and B(106)) xor (A(39) and B(105)) xor (A(40) and B(104)) xor (A(41) and B(103)) xor (A(42) and B(102)) xor (A(43) and B(101)) xor (A(44) and B(100)) xor (A(45) and B(99)) xor (A(46) and B(98)) xor (A(47) and B(97)) xor (A(48) and B(96)) xor (A(49) and B(95)) xor (A(50) and B(94)) xor (A(51) and B(93)) xor (A(52) and B(92)) xor (A(53) and B(91)) xor (A(54) and B(90)) xor (A(55) and B(89)) xor (A(56) and B(88)) xor (A(57) and B(87)) xor (A(58) and B(86)) xor (A(59) and B(85)) xor (A(60) and B(84)) xor (A(61) and B(83)) xor (A(62) and B(82)) xor (A(63) and B(81)) xor (A(64) and B(80)) xor (A(65) and B(79)) xor (A(66) and B(78)) xor (A(67) and B(77)) xor (A(68) and B(76)) xor (A(69) and B(75)) xor (A(70) and B(74)) xor (A(71) and B(73)) xor (A(72) and B(72)) xor (A(73) and B(71)) xor (A(74) and B(70)) xor (A(75) and B(69)) xor (A(76) and B(68)) xor (A(77) and B(67)) xor (A(78) and B(66)) xor (A(79) and B(65)) xor (A(80) and B(64)) xor (A(81) and B(63)) xor (A(82) and B(62)) xor (A(83) and B(61)) xor (A(84) and B(60)) xor (A(85) and B(59)) xor (A(86) and B(58)) xor (A(87) and B(57)) xor (A(88) and B(56)) xor (A(89) and B(55)) xor (A(90) and B(54)) xor (A(91) and B(53)) xor (A(92) and B(52)) xor (A(93) and B(51)) xor (A(94) and B(50)) xor (A(95) and B(49)) xor (A(96) and B(48)) xor (A(97) and B(47)) xor (A(98) and B(46)) xor (A(99) and B(45)) xor (A(100) and B(44)) xor (A(101) and B(43)) xor (A(102) and B(42)) xor (A(103) and B(41)) xor (A(104) and B(40)) xor (A(105) and B(39)) xor (A(106) and B(38)) xor (A(107) and B(37)) xor (A(108) and B(36)) xor (A(109) and B(35)) xor (A(110) and B(34)) xor (A(111) and B(33)) xor (A(112) and B(32)) xor (A(113) and B(31)) xor (A(114) and B(30)) xor (A(115) and B(29)) xor (A(116) and B(28)) xor (A(117) and B(27)) xor (A(118) and B(26)) xor (A(119) and B(25)) xor (A(120) and B(24)) xor (A(121) and B(23)) xor (A(122) and B(23)) xor (A(123) and B(21)) xor (A(124) and B(20)) xor (A(125) and B(19)) xor (A(126) and B(18)) xor (A(23) and B(127)) xor (A(23) and B(126)) xor (A(24) and B(125)) xor (A(25) and B(124)) xor (A(26) and B(123)) xor (A(27) and B(122)) xor (A(28) and B(121)) xor (A(29) and B(120)) xor (A(30) and B(119)) xor (A(31) and B(118)) xor (A(32) and B(117)) xor (A(33) and B(116)) xor (A(34) and B(115)) xor (A(35) and B(114)) xor (A(36) and B(113)) xor (A(37) and B(112)) xor (A(38) and B(111)) xor (A(39) and B(110)) xor (A(40) and B(109)) xor (A(41) and B(108)) xor (A(42) and B(107)) xor (A(43) and B(106)) xor (A(44) and B(105)) xor (A(45) and B(104)) xor (A(46) and B(103)) xor (A(47) and B(102)) xor (A(48) and B(101)) xor (A(49) and B(100)) xor (A(50) and B(99)) xor (A(51) and B(98)) xor (A(52) and B(97)) xor (A(53) and B(96)) xor (A(54) and B(95)) xor (A(55) and B(94)) xor (A(56) and B(93)) xor (A(57) and B(92)) xor (A(58) and B(91)) xor (A(59) and B(90)) xor (A(60) and B(89)) xor (A(61) and B(88)) xor (A(62) and B(87)) xor (A(63) and B(86)) xor (A(64) and B(85)) xor (A(65) and B(84)) xor (A(66) and B(83)) xor (A(67) and B(82)) xor (A(68) and B(81)) xor (A(69) and B(80)) xor (A(70) and B(79)) xor (A(71) and B(78)) xor (A(72) and B(77)) xor (A(73) and B(76)) xor (A(74) and B(75)) xor (A(75) and B(74)) xor (A(76) and B(73)) xor (A(77) and B(72)) xor (A(78) and B(71)) xor (A(79) and B(70)) xor (A(80) and B(69)) xor (A(81) and B(68)) xor (A(82) and B(67)) xor (A(83) and B(66)) xor (A(84) and B(65)) xor (A(85) and B(64)) xor (A(86) and B(63)) xor (A(87) and B(62)) xor (A(88) and B(61)) xor (A(89) and B(60)) xor (A(90) and B(59)) xor (A(91) and B(58)) xor (A(92) and B(57)) xor (A(93) and B(56)) xor (A(94) and B(55)) xor (A(95) and B(54)) xor (A(96) and B(53)) xor (A(97) and B(52)) xor (A(98) and B(51)) xor (A(99) and B(50)) xor (A(100) and B(49)) xor (A(101) and B(48)) xor (A(102) and B(47)) xor (A(103) and B(46)) xor (A(104) and B(45)) xor (A(105) and B(44)) xor (A(106) and B(43)) xor (A(107) and B(42)) xor (A(108) and B(41)) xor (A(109) and B(40)) xor (A(110) and B(39)) xor (A(111) and B(38)) xor (A(112) and B(37)) xor (A(113) and B(36)) xor (A(114) and B(35)) xor (A(115) and B(34)) xor (A(116) and B(33)) xor (A(117) and B(32)) xor (A(118) and B(31)) xor (A(119) and B(30)) xor (A(120) and B(29)) xor (A(121) and B(28)) xor (A(122) and B(27)) xor (A(123) and B(26)) xor (A(124) and B(25)) xor (A(125) and B(24)) xor (A(126) and B(23)) xor (A(23) and B(127)) xor (A(24) and B(126)) xor (A(25) and B(125)) xor (A(26) and B(124)) xor (A(27) and B(123)) xor (A(28) and B(122)) xor (A(29) and B(121)) xor (A(30) and B(120)) xor (A(31) and B(119)) xor (A(32) and B(118)) xor (A(33) and B(117)) xor (A(34) and B(116)) xor (A(35) and B(115)) xor (A(36) and B(114)) xor (A(37) and B(113)) xor (A(38) and B(112)) xor (A(39) and B(111)) xor (A(40) and B(110)) xor (A(41) and B(109)) xor (A(42) and B(108)) xor (A(43) and B(107)) xor (A(44) and B(106)) xor (A(45) and B(105)) xor (A(46) and B(104)) xor (A(47) and B(103)) xor (A(48) and B(102)) xor (A(49) and B(101)) xor (A(50) and B(100)) xor (A(51) and B(99)) xor (A(52) and B(98)) xor (A(53) and B(97)) xor (A(54) and B(96)) xor (A(55) and B(95)) xor (A(56) and B(94)) xor (A(57) and B(93)) xor (A(58) and B(92)) xor (A(59) and B(91)) xor (A(60) and B(90)) xor (A(61) and B(89)) xor (A(62) and B(88)) xor (A(63) and B(87)) xor (A(64) and B(86)) xor (A(65) and B(85)) xor (A(66) and B(84)) xor (A(67) and B(83)) xor (A(68) and B(82)) xor (A(69) and B(81)) xor (A(70) and B(80)) xor (A(71) and B(79)) xor (A(72) and B(78)) xor (A(73) and B(77)) xor (A(74) and B(76)) xor (A(75) and B(75)) xor (A(76) and B(74)) xor (A(77) and B(73)) xor (A(78) and B(72)) xor (A(79) and B(71)) xor (A(80) and B(70)) xor (A(81) and B(69)) xor (A(82) and B(68)) xor (A(83) and B(67)) xor (A(84) and B(66)) xor (A(85) and B(65)) xor (A(86) and B(64)) xor (A(87) and B(63)) xor (A(88) and B(62)) xor (A(89) and B(61)) xor (A(90) and B(60)) xor (A(91) and B(59)) xor (A(92) and B(58)) xor (A(93) and B(57)) xor (A(94) and B(56)) xor (A(95) and B(55)) xor (A(96) and B(54)) xor (A(97) and B(53)) xor (A(98) and B(52)) xor (A(99) and B(51)) xor (A(100) and B(50)) xor (A(101) and B(49)) xor (A(102) and B(48)) xor (A(103) and B(47)) xor (A(104) and B(46)) xor (A(105) and B(45)) xor (A(106) and B(44)) xor (A(107) and B(43)) xor (A(108) and B(42)) xor (A(109) and B(41)) xor (A(110) and B(40)) xor (A(111) and B(39)) xor (A(112) and B(38)) xor (A(113) and B(37)) xor (A(114) and B(36)) xor (A(115) and B(35)) xor (A(116) and B(34)) xor (A(117) and B(33)) xor (A(118) and B(32)) xor (A(119) and B(31)) xor (A(120) and B(30)) xor (A(121) and B(29)) xor (A(122) and B(28)) xor (A(123) and B(27)) xor (A(124) and B(26)) xor (A(125) and B(25)) xor (A(126) and B(24)) xor (A(24) and B(127)) xor (A(25) and B(126)) xor (A(26) and B(125)) xor (A(27) and B(124)) xor (A(28) and B(123)) xor (A(29) and B(122)) xor (A(30) and B(121)) xor (A(31) and B(120)) xor (A(32) and B(119)) xor (A(33) and B(118)) xor (A(34) and B(117)) xor (A(35) and B(116)) xor (A(36) and B(115)) xor (A(37) and B(114)) xor (A(38) and B(113)) xor (A(39) and B(112)) xor (A(40) and B(111)) xor (A(41) and B(110)) xor (A(42) and B(109)) xor (A(43) and B(108)) xor (A(44) and B(107)) xor (A(45) and B(106)) xor (A(46) and B(105)) xor (A(47) and B(104)) xor (A(48) and B(103)) xor (A(49) and B(102)) xor (A(50) and B(101)) xor (A(51) and B(100)) xor (A(52) and B(99)) xor (A(53) and B(98)) xor (A(54) and B(97)) xor (A(55) and B(96)) xor (A(56) and B(95)) xor (A(57) and B(94)) xor (A(58) and B(93)) xor (A(59) and B(92)) xor (A(60) and B(91)) xor (A(61) and B(90)) xor (A(62) and B(89)) xor (A(63) and B(88)) xor (A(64) and B(87)) xor (A(65) and B(86)) xor (A(66) and B(85)) xor (A(67) and B(84)) xor (A(68) and B(83)) xor (A(69) and B(82)) xor (A(70) and B(81)) xor (A(71) and B(80)) xor (A(72) and B(79)) xor (A(73) and B(78)) xor (A(74) and B(77)) xor (A(75) and B(76)) xor (A(76) and B(75)) xor (A(77) and B(74)) xor (A(78) and B(73)) xor (A(79) and B(72)) xor (A(80) and B(71)) xor (A(81) and B(70)) xor (A(82) and B(69)) xor (A(83) and B(68)) xor (A(84) and B(67)) xor (A(85) and B(66)) xor (A(86) and B(65)) xor (A(87) and B(64)) xor (A(88) and B(63)) xor (A(89) and B(62)) xor (A(90) and B(61)) xor (A(91) and B(60)) xor (A(92) and B(59)) xor (A(93) and B(58)) xor (A(94) and B(57)) xor (A(95) and B(56)) xor (A(96) and B(55)) xor (A(97) and B(54)) xor (A(98) and B(53)) xor (A(99) and B(52)) xor (A(100) and B(51)) xor (A(101) and B(50)) xor (A(102) and B(49)) xor (A(103) and B(48)) xor (A(104) and B(47)) xor (A(105) and B(46)) xor (A(106) and B(45)) xor (A(107) and B(44)) xor (A(108) and B(43)) xor (A(109) and B(42)) xor (A(110) and B(41)) xor (A(111) and B(40)) xor (A(112) and B(39)) xor (A(113) and B(38)) xor (A(114) and B(37)) xor (A(115) and B(36)) xor (A(116) and B(35)) xor (A(117) and B(34)) xor (A(118) and B(33)) xor (A(119) and B(32)) xor (A(120) and B(31)) xor (A(121) and B(30)) xor (A(122) and B(29)) xor (A(123) and B(28)) xor (A(124) and B(27)) xor (A(125) and B(26)) xor (A(126) and B(26));
    C(25)  <= (A(0) and B(25)) xor (A(1) and B(24)) xor (A(2) and B(23)) xor (A(3) and B(23)) xor (A(4) and B(21)) xor (A(5) and B(20)) xor (A(6) and B(19)) xor (A(7) and B(18)) xor (A(8) and B(17)) xor (A(9) and B(16)) xor (A(10) and B(15)) xor (A(11) and B(14)) xor (A(12) and B(13)) xor (A(13) and B(12)) xor (A(14) and B(11)) xor (A(15) and B(10)) xor (A(16) and B(9)) xor (A(17) and B(8)) xor (A(18) and B(7)) xor (A(19) and B(6)) xor (A(20) and B(5)) xor (A(21) and B(4)) xor (A(23) and B(3)) xor (A(23) and B(2)) xor (A(24) and B(1)) xor (A(25) and B(0)) xor (A(18) and B(127)) xor (A(19) and B(126)) xor (A(20) and B(125)) xor (A(21) and B(124)) xor (A(23) and B(123)) xor (A(23) and B(122)) xor (A(24) and B(121)) xor (A(25) and B(120)) xor (A(26) and B(119)) xor (A(27) and B(118)) xor (A(28) and B(117)) xor (A(29) and B(116)) xor (A(30) and B(115)) xor (A(31) and B(114)) xor (A(32) and B(113)) xor (A(33) and B(112)) xor (A(34) and B(111)) xor (A(35) and B(110)) xor (A(36) and B(109)) xor (A(37) and B(108)) xor (A(38) and B(107)) xor (A(39) and B(106)) xor (A(40) and B(105)) xor (A(41) and B(104)) xor (A(42) and B(103)) xor (A(43) and B(102)) xor (A(44) and B(101)) xor (A(45) and B(100)) xor (A(46) and B(99)) xor (A(47) and B(98)) xor (A(48) and B(97)) xor (A(49) and B(96)) xor (A(50) and B(95)) xor (A(51) and B(94)) xor (A(52) and B(93)) xor (A(53) and B(92)) xor (A(54) and B(91)) xor (A(55) and B(90)) xor (A(56) and B(89)) xor (A(57) and B(88)) xor (A(58) and B(87)) xor (A(59) and B(86)) xor (A(60) and B(85)) xor (A(61) and B(84)) xor (A(62) and B(83)) xor (A(63) and B(82)) xor (A(64) and B(81)) xor (A(65) and B(80)) xor (A(66) and B(79)) xor (A(67) and B(78)) xor (A(68) and B(77)) xor (A(69) and B(76)) xor (A(70) and B(75)) xor (A(71) and B(74)) xor (A(72) and B(73)) xor (A(73) and B(72)) xor (A(74) and B(71)) xor (A(75) and B(70)) xor (A(76) and B(69)) xor (A(77) and B(68)) xor (A(78) and B(67)) xor (A(79) and B(66)) xor (A(80) and B(65)) xor (A(81) and B(64)) xor (A(82) and B(63)) xor (A(83) and B(62)) xor (A(84) and B(61)) xor (A(85) and B(60)) xor (A(86) and B(59)) xor (A(87) and B(58)) xor (A(88) and B(57)) xor (A(89) and B(56)) xor (A(90) and B(55)) xor (A(91) and B(54)) xor (A(92) and B(53)) xor (A(93) and B(52)) xor (A(94) and B(51)) xor (A(95) and B(50)) xor (A(96) and B(49)) xor (A(97) and B(48)) xor (A(98) and B(47)) xor (A(99) and B(46)) xor (A(100) and B(45)) xor (A(101) and B(44)) xor (A(102) and B(43)) xor (A(103) and B(42)) xor (A(104) and B(41)) xor (A(105) and B(40)) xor (A(106) and B(39)) xor (A(107) and B(38)) xor (A(108) and B(37)) xor (A(109) and B(36)) xor (A(110) and B(35)) xor (A(111) and B(34)) xor (A(112) and B(33)) xor (A(113) and B(32)) xor (A(114) and B(31)) xor (A(115) and B(30)) xor (A(116) and B(29)) xor (A(117) and B(28)) xor (A(118) and B(27)) xor (A(119) and B(26)) xor (A(120) and B(25)) xor (A(121) and B(24)) xor (A(122) and B(23)) xor (A(123) and B(23)) xor (A(124) and B(21)) xor (A(125) and B(20)) xor (A(126) and B(19)) xor (A(23) and B(127)) xor (A(24) and B(126)) xor (A(25) and B(125)) xor (A(26) and B(124)) xor (A(27) and B(123)) xor (A(28) and B(122)) xor (A(29) and B(121)) xor (A(30) and B(120)) xor (A(31) and B(119)) xor (A(32) and B(118)) xor (A(33) and B(117)) xor (A(34) and B(116)) xor (A(35) and B(115)) xor (A(36) and B(114)) xor (A(37) and B(113)) xor (A(38) and B(112)) xor (A(39) and B(111)) xor (A(40) and B(110)) xor (A(41) and B(109)) xor (A(42) and B(108)) xor (A(43) and B(107)) xor (A(44) and B(106)) xor (A(45) and B(105)) xor (A(46) and B(104)) xor (A(47) and B(103)) xor (A(48) and B(102)) xor (A(49) and B(101)) xor (A(50) and B(100)) xor (A(51) and B(99)) xor (A(52) and B(98)) xor (A(53) and B(97)) xor (A(54) and B(96)) xor (A(55) and B(95)) xor (A(56) and B(94)) xor (A(57) and B(93)) xor (A(58) and B(92)) xor (A(59) and B(91)) xor (A(60) and B(90)) xor (A(61) and B(89)) xor (A(62) and B(88)) xor (A(63) and B(87)) xor (A(64) and B(86)) xor (A(65) and B(85)) xor (A(66) and B(84)) xor (A(67) and B(83)) xor (A(68) and B(82)) xor (A(69) and B(81)) xor (A(70) and B(80)) xor (A(71) and B(79)) xor (A(72) and B(78)) xor (A(73) and B(77)) xor (A(74) and B(76)) xor (A(75) and B(75)) xor (A(76) and B(74)) xor (A(77) and B(73)) xor (A(78) and B(72)) xor (A(79) and B(71)) xor (A(80) and B(70)) xor (A(81) and B(69)) xor (A(82) and B(68)) xor (A(83) and B(67)) xor (A(84) and B(66)) xor (A(85) and B(65)) xor (A(86) and B(64)) xor (A(87) and B(63)) xor (A(88) and B(62)) xor (A(89) and B(61)) xor (A(90) and B(60)) xor (A(91) and B(59)) xor (A(92) and B(58)) xor (A(93) and B(57)) xor (A(94) and B(56)) xor (A(95) and B(55)) xor (A(96) and B(54)) xor (A(97) and B(53)) xor (A(98) and B(52)) xor (A(99) and B(51)) xor (A(100) and B(50)) xor (A(101) and B(49)) xor (A(102) and B(48)) xor (A(103) and B(47)) xor (A(104) and B(46)) xor (A(105) and B(45)) xor (A(106) and B(44)) xor (A(107) and B(43)) xor (A(108) and B(42)) xor (A(109) and B(41)) xor (A(110) and B(40)) xor (A(111) and B(39)) xor (A(112) and B(38)) xor (A(113) and B(37)) xor (A(114) and B(36)) xor (A(115) and B(35)) xor (A(116) and B(34)) xor (A(117) and B(33)) xor (A(118) and B(32)) xor (A(119) and B(31)) xor (A(120) and B(30)) xor (A(121) and B(29)) xor (A(122) and B(28)) xor (A(123) and B(27)) xor (A(124) and B(26)) xor (A(125) and B(25)) xor (A(126) and B(24)) xor (A(24) and B(127)) xor (A(25) and B(126)) xor (A(26) and B(125)) xor (A(27) and B(124)) xor (A(28) and B(123)) xor (A(29) and B(122)) xor (A(30) and B(121)) xor (A(31) and B(120)) xor (A(32) and B(119)) xor (A(33) and B(118)) xor (A(34) and B(117)) xor (A(35) and B(116)) xor (A(36) and B(115)) xor (A(37) and B(114)) xor (A(38) and B(113)) xor (A(39) and B(112)) xor (A(40) and B(111)) xor (A(41) and B(110)) xor (A(42) and B(109)) xor (A(43) and B(108)) xor (A(44) and B(107)) xor (A(45) and B(106)) xor (A(46) and B(105)) xor (A(47) and B(104)) xor (A(48) and B(103)) xor (A(49) and B(102)) xor (A(50) and B(101)) xor (A(51) and B(100)) xor (A(52) and B(99)) xor (A(53) and B(98)) xor (A(54) and B(97)) xor (A(55) and B(96)) xor (A(56) and B(95)) xor (A(57) and B(94)) xor (A(58) and B(93)) xor (A(59) and B(92)) xor (A(60) and B(91)) xor (A(61) and B(90)) xor (A(62) and B(89)) xor (A(63) and B(88)) xor (A(64) and B(87)) xor (A(65) and B(86)) xor (A(66) and B(85)) xor (A(67) and B(84)) xor (A(68) and B(83)) xor (A(69) and B(82)) xor (A(70) and B(81)) xor (A(71) and B(80)) xor (A(72) and B(79)) xor (A(73) and B(78)) xor (A(74) and B(77)) xor (A(75) and B(76)) xor (A(76) and B(75)) xor (A(77) and B(74)) xor (A(78) and B(73)) xor (A(79) and B(72)) xor (A(80) and B(71)) xor (A(81) and B(70)) xor (A(82) and B(69)) xor (A(83) and B(68)) xor (A(84) and B(67)) xor (A(85) and B(66)) xor (A(86) and B(65)) xor (A(87) and B(64)) xor (A(88) and B(63)) xor (A(89) and B(62)) xor (A(90) and B(61)) xor (A(91) and B(60)) xor (A(92) and B(59)) xor (A(93) and B(58)) xor (A(94) and B(57)) xor (A(95) and B(56)) xor (A(96) and B(55)) xor (A(97) and B(54)) xor (A(98) and B(53)) xor (A(99) and B(52)) xor (A(100) and B(51)) xor (A(101) and B(50)) xor (A(102) and B(49)) xor (A(103) and B(48)) xor (A(104) and B(47)) xor (A(105) and B(46)) xor (A(106) and B(45)) xor (A(107) and B(44)) xor (A(108) and B(43)) xor (A(109) and B(42)) xor (A(110) and B(41)) xor (A(111) and B(40)) xor (A(112) and B(39)) xor (A(113) and B(38)) xor (A(114) and B(37)) xor (A(115) and B(36)) xor (A(116) and B(35)) xor (A(117) and B(34)) xor (A(118) and B(33)) xor (A(119) and B(32)) xor (A(120) and B(31)) xor (A(121) and B(30)) xor (A(122) and B(29)) xor (A(123) and B(28)) xor (A(124) and B(27)) xor (A(125) and B(26)) xor (A(126) and B(25)) xor (A(25) and B(127)) xor (A(26) and B(126)) xor (A(27) and B(125)) xor (A(28) and B(124)) xor (A(29) and B(123)) xor (A(30) and B(122)) xor (A(31) and B(121)) xor (A(32) and B(120)) xor (A(33) and B(119)) xor (A(34) and B(118)) xor (A(35) and B(117)) xor (A(36) and B(116)) xor (A(37) and B(115)) xor (A(38) and B(114)) xor (A(39) and B(113)) xor (A(40) and B(112)) xor (A(41) and B(111)) xor (A(42) and B(110)) xor (A(43) and B(109)) xor (A(44) and B(108)) xor (A(45) and B(107)) xor (A(46) and B(106)) xor (A(47) and B(105)) xor (A(48) and B(104)) xor (A(49) and B(103)) xor (A(50) and B(102)) xor (A(51) and B(101)) xor (A(52) and B(100)) xor (A(53) and B(99)) xor (A(54) and B(98)) xor (A(55) and B(97)) xor (A(56) and B(96)) xor (A(57) and B(95)) xor (A(58) and B(94)) xor (A(59) and B(93)) xor (A(60) and B(92)) xor (A(61) and B(91)) xor (A(62) and B(90)) xor (A(63) and B(89)) xor (A(64) and B(88)) xor (A(65) and B(87)) xor (A(66) and B(86)) xor (A(67) and B(85)) xor (A(68) and B(84)) xor (A(69) and B(83)) xor (A(70) and B(82)) xor (A(71) and B(81)) xor (A(72) and B(80)) xor (A(73) and B(79)) xor (A(74) and B(78)) xor (A(75) and B(77)) xor (A(76) and B(76)) xor (A(77) and B(75)) xor (A(78) and B(74)) xor (A(79) and B(73)) xor (A(80) and B(72)) xor (A(81) and B(71)) xor (A(82) and B(70)) xor (A(83) and B(69)) xor (A(84) and B(68)) xor (A(85) and B(67)) xor (A(86) and B(66)) xor (A(87) and B(65)) xor (A(88) and B(64)) xor (A(89) and B(63)) xor (A(90) and B(62)) xor (A(91) and B(61)) xor (A(92) and B(60)) xor (A(93) and B(59)) xor (A(94) and B(58)) xor (A(95) and B(57)) xor (A(96) and B(56)) xor (A(97) and B(55)) xor (A(98) and B(54)) xor (A(99) and B(53)) xor (A(100) and B(52)) xor (A(101) and B(51)) xor (A(102) and B(50)) xor (A(103) and B(49)) xor (A(104) and B(48)) xor (A(105) and B(47)) xor (A(106) and B(46)) xor (A(107) and B(45)) xor (A(108) and B(44)) xor (A(109) and B(43)) xor (A(110) and B(42)) xor (A(111) and B(41)) xor (A(112) and B(40)) xor (A(113) and B(39)) xor (A(114) and B(38)) xor (A(115) and B(37)) xor (A(116) and B(36)) xor (A(117) and B(35)) xor (A(118) and B(34)) xor (A(119) and B(33)) xor (A(120) and B(32)) xor (A(121) and B(31)) xor (A(122) and B(30)) xor (A(123) and B(29)) xor (A(124) and B(28)) xor (A(125) and B(27)) xor (A(126) and B(27));
    C(26)  <= (A(0) and B(26)) xor (A(1) and B(25)) xor (A(2) and B(24)) xor (A(3) and B(23)) xor (A(4) and B(23)) xor (A(5) and B(21)) xor (A(6) and B(20)) xor (A(7) and B(19)) xor (A(8) and B(18)) xor (A(9) and B(17)) xor (A(10) and B(16)) xor (A(11) and B(15)) xor (A(12) and B(14)) xor (A(13) and B(13)) xor (A(14) and B(12)) xor (A(15) and B(11)) xor (A(16) and B(10)) xor (A(17) and B(9)) xor (A(18) and B(8)) xor (A(19) and B(7)) xor (A(20) and B(6)) xor (A(21) and B(5)) xor (A(23) and B(4)) xor (A(23) and B(3)) xor (A(24) and B(2)) xor (A(25) and B(1)) xor (A(26) and B(0)) xor (A(19) and B(127)) xor (A(20) and B(126)) xor (A(21) and B(125)) xor (A(23) and B(124)) xor (A(23) and B(123)) xor (A(24) and B(122)) xor (A(25) and B(121)) xor (A(26) and B(120)) xor (A(27) and B(119)) xor (A(28) and B(118)) xor (A(29) and B(117)) xor (A(30) and B(116)) xor (A(31) and B(115)) xor (A(32) and B(114)) xor (A(33) and B(113)) xor (A(34) and B(112)) xor (A(35) and B(111)) xor (A(36) and B(110)) xor (A(37) and B(109)) xor (A(38) and B(108)) xor (A(39) and B(107)) xor (A(40) and B(106)) xor (A(41) and B(105)) xor (A(42) and B(104)) xor (A(43) and B(103)) xor (A(44) and B(102)) xor (A(45) and B(101)) xor (A(46) and B(100)) xor (A(47) and B(99)) xor (A(48) and B(98)) xor (A(49) and B(97)) xor (A(50) and B(96)) xor (A(51) and B(95)) xor (A(52) and B(94)) xor (A(53) and B(93)) xor (A(54) and B(92)) xor (A(55) and B(91)) xor (A(56) and B(90)) xor (A(57) and B(89)) xor (A(58) and B(88)) xor (A(59) and B(87)) xor (A(60) and B(86)) xor (A(61) and B(85)) xor (A(62) and B(84)) xor (A(63) and B(83)) xor (A(64) and B(82)) xor (A(65) and B(81)) xor (A(66) and B(80)) xor (A(67) and B(79)) xor (A(68) and B(78)) xor (A(69) and B(77)) xor (A(70) and B(76)) xor (A(71) and B(75)) xor (A(72) and B(74)) xor (A(73) and B(73)) xor (A(74) and B(72)) xor (A(75) and B(71)) xor (A(76) and B(70)) xor (A(77) and B(69)) xor (A(78) and B(68)) xor (A(79) and B(67)) xor (A(80) and B(66)) xor (A(81) and B(65)) xor (A(82) and B(64)) xor (A(83) and B(63)) xor (A(84) and B(62)) xor (A(85) and B(61)) xor (A(86) and B(60)) xor (A(87) and B(59)) xor (A(88) and B(58)) xor (A(89) and B(57)) xor (A(90) and B(56)) xor (A(91) and B(55)) xor (A(92) and B(54)) xor (A(93) and B(53)) xor (A(94) and B(52)) xor (A(95) and B(51)) xor (A(96) and B(50)) xor (A(97) and B(49)) xor (A(98) and B(48)) xor (A(99) and B(47)) xor (A(100) and B(46)) xor (A(101) and B(45)) xor (A(102) and B(44)) xor (A(103) and B(43)) xor (A(104) and B(42)) xor (A(105) and B(41)) xor (A(106) and B(40)) xor (A(107) and B(39)) xor (A(108) and B(38)) xor (A(109) and B(37)) xor (A(110) and B(36)) xor (A(111) and B(35)) xor (A(112) and B(34)) xor (A(113) and B(33)) xor (A(114) and B(32)) xor (A(115) and B(31)) xor (A(116) and B(30)) xor (A(117) and B(29)) xor (A(118) and B(28)) xor (A(119) and B(27)) xor (A(120) and B(26)) xor (A(121) and B(25)) xor (A(122) and B(24)) xor (A(123) and B(23)) xor (A(124) and B(23)) xor (A(125) and B(21)) xor (A(126) and B(20)) xor (A(24) and B(127)) xor (A(25) and B(126)) xor (A(26) and B(125)) xor (A(27) and B(124)) xor (A(28) and B(123)) xor (A(29) and B(122)) xor (A(30) and B(121)) xor (A(31) and B(120)) xor (A(32) and B(119)) xor (A(33) and B(118)) xor (A(34) and B(117)) xor (A(35) and B(116)) xor (A(36) and B(115)) xor (A(37) and B(114)) xor (A(38) and B(113)) xor (A(39) and B(112)) xor (A(40) and B(111)) xor (A(41) and B(110)) xor (A(42) and B(109)) xor (A(43) and B(108)) xor (A(44) and B(107)) xor (A(45) and B(106)) xor (A(46) and B(105)) xor (A(47) and B(104)) xor (A(48) and B(103)) xor (A(49) and B(102)) xor (A(50) and B(101)) xor (A(51) and B(100)) xor (A(52) and B(99)) xor (A(53) and B(98)) xor (A(54) and B(97)) xor (A(55) and B(96)) xor (A(56) and B(95)) xor (A(57) and B(94)) xor (A(58) and B(93)) xor (A(59) and B(92)) xor (A(60) and B(91)) xor (A(61) and B(90)) xor (A(62) and B(89)) xor (A(63) and B(88)) xor (A(64) and B(87)) xor (A(65) and B(86)) xor (A(66) and B(85)) xor (A(67) and B(84)) xor (A(68) and B(83)) xor (A(69) and B(82)) xor (A(70) and B(81)) xor (A(71) and B(80)) xor (A(72) and B(79)) xor (A(73) and B(78)) xor (A(74) and B(77)) xor (A(75) and B(76)) xor (A(76) and B(75)) xor (A(77) and B(74)) xor (A(78) and B(73)) xor (A(79) and B(72)) xor (A(80) and B(71)) xor (A(81) and B(70)) xor (A(82) and B(69)) xor (A(83) and B(68)) xor (A(84) and B(67)) xor (A(85) and B(66)) xor (A(86) and B(65)) xor (A(87) and B(64)) xor (A(88) and B(63)) xor (A(89) and B(62)) xor (A(90) and B(61)) xor (A(91) and B(60)) xor (A(92) and B(59)) xor (A(93) and B(58)) xor (A(94) and B(57)) xor (A(95) and B(56)) xor (A(96) and B(55)) xor (A(97) and B(54)) xor (A(98) and B(53)) xor (A(99) and B(52)) xor (A(100) and B(51)) xor (A(101) and B(50)) xor (A(102) and B(49)) xor (A(103) and B(48)) xor (A(104) and B(47)) xor (A(105) and B(46)) xor (A(106) and B(45)) xor (A(107) and B(44)) xor (A(108) and B(43)) xor (A(109) and B(42)) xor (A(110) and B(41)) xor (A(111) and B(40)) xor (A(112) and B(39)) xor (A(113) and B(38)) xor (A(114) and B(37)) xor (A(115) and B(36)) xor (A(116) and B(35)) xor (A(117) and B(34)) xor (A(118) and B(33)) xor (A(119) and B(32)) xor (A(120) and B(31)) xor (A(121) and B(30)) xor (A(122) and B(29)) xor (A(123) and B(28)) xor (A(124) and B(27)) xor (A(125) and B(26)) xor (A(126) and B(25)) xor (A(25) and B(127)) xor (A(26) and B(126)) xor (A(27) and B(125)) xor (A(28) and B(124)) xor (A(29) and B(123)) xor (A(30) and B(122)) xor (A(31) and B(121)) xor (A(32) and B(120)) xor (A(33) and B(119)) xor (A(34) and B(118)) xor (A(35) and B(117)) xor (A(36) and B(116)) xor (A(37) and B(115)) xor (A(38) and B(114)) xor (A(39) and B(113)) xor (A(40) and B(112)) xor (A(41) and B(111)) xor (A(42) and B(110)) xor (A(43) and B(109)) xor (A(44) and B(108)) xor (A(45) and B(107)) xor (A(46) and B(106)) xor (A(47) and B(105)) xor (A(48) and B(104)) xor (A(49) and B(103)) xor (A(50) and B(102)) xor (A(51) and B(101)) xor (A(52) and B(100)) xor (A(53) and B(99)) xor (A(54) and B(98)) xor (A(55) and B(97)) xor (A(56) and B(96)) xor (A(57) and B(95)) xor (A(58) and B(94)) xor (A(59) and B(93)) xor (A(60) and B(92)) xor (A(61) and B(91)) xor (A(62) and B(90)) xor (A(63) and B(89)) xor (A(64) and B(88)) xor (A(65) and B(87)) xor (A(66) and B(86)) xor (A(67) and B(85)) xor (A(68) and B(84)) xor (A(69) and B(83)) xor (A(70) and B(82)) xor (A(71) and B(81)) xor (A(72) and B(80)) xor (A(73) and B(79)) xor (A(74) and B(78)) xor (A(75) and B(77)) xor (A(76) and B(76)) xor (A(77) and B(75)) xor (A(78) and B(74)) xor (A(79) and B(73)) xor (A(80) and B(72)) xor (A(81) and B(71)) xor (A(82) and B(70)) xor (A(83) and B(69)) xor (A(84) and B(68)) xor (A(85) and B(67)) xor (A(86) and B(66)) xor (A(87) and B(65)) xor (A(88) and B(64)) xor (A(89) and B(63)) xor (A(90) and B(62)) xor (A(91) and B(61)) xor (A(92) and B(60)) xor (A(93) and B(59)) xor (A(94) and B(58)) xor (A(95) and B(57)) xor (A(96) and B(56)) xor (A(97) and B(55)) xor (A(98) and B(54)) xor (A(99) and B(53)) xor (A(100) and B(52)) xor (A(101) and B(51)) xor (A(102) and B(50)) xor (A(103) and B(49)) xor (A(104) and B(48)) xor (A(105) and B(47)) xor (A(106) and B(46)) xor (A(107) and B(45)) xor (A(108) and B(44)) xor (A(109) and B(43)) xor (A(110) and B(42)) xor (A(111) and B(41)) xor (A(112) and B(40)) xor (A(113) and B(39)) xor (A(114) and B(38)) xor (A(115) and B(37)) xor (A(116) and B(36)) xor (A(117) and B(35)) xor (A(118) and B(34)) xor (A(119) and B(33)) xor (A(120) and B(32)) xor (A(121) and B(31)) xor (A(122) and B(30)) xor (A(123) and B(29)) xor (A(124) and B(28)) xor (A(125) and B(27)) xor (A(126) and B(26)) xor (A(26) and B(127)) xor (A(27) and B(126)) xor (A(28) and B(125)) xor (A(29) and B(124)) xor (A(30) and B(123)) xor (A(31) and B(122)) xor (A(32) and B(121)) xor (A(33) and B(120)) xor (A(34) and B(119)) xor (A(35) and B(118)) xor (A(36) and B(117)) xor (A(37) and B(116)) xor (A(38) and B(115)) xor (A(39) and B(114)) xor (A(40) and B(113)) xor (A(41) and B(112)) xor (A(42) and B(111)) xor (A(43) and B(110)) xor (A(44) and B(109)) xor (A(45) and B(108)) xor (A(46) and B(107)) xor (A(47) and B(106)) xor (A(48) and B(105)) xor (A(49) and B(104)) xor (A(50) and B(103)) xor (A(51) and B(102)) xor (A(52) and B(101)) xor (A(53) and B(100)) xor (A(54) and B(99)) xor (A(55) and B(98)) xor (A(56) and B(97)) xor (A(57) and B(96)) xor (A(58) and B(95)) xor (A(59) and B(94)) xor (A(60) and B(93)) xor (A(61) and B(92)) xor (A(62) and B(91)) xor (A(63) and B(90)) xor (A(64) and B(89)) xor (A(65) and B(88)) xor (A(66) and B(87)) xor (A(67) and B(86)) xor (A(68) and B(85)) xor (A(69) and B(84)) xor (A(70) and B(83)) xor (A(71) and B(82)) xor (A(72) and B(81)) xor (A(73) and B(80)) xor (A(74) and B(79)) xor (A(75) and B(78)) xor (A(76) and B(77)) xor (A(77) and B(76)) xor (A(78) and B(75)) xor (A(79) and B(74)) xor (A(80) and B(73)) xor (A(81) and B(72)) xor (A(82) and B(71)) xor (A(83) and B(70)) xor (A(84) and B(69)) xor (A(85) and B(68)) xor (A(86) and B(67)) xor (A(87) and B(66)) xor (A(88) and B(65)) xor (A(89) and B(64)) xor (A(90) and B(63)) xor (A(91) and B(62)) xor (A(92) and B(61)) xor (A(93) and B(60)) xor (A(94) and B(59)) xor (A(95) and B(58)) xor (A(96) and B(57)) xor (A(97) and B(56)) xor (A(98) and B(55)) xor (A(99) and B(54)) xor (A(100) and B(53)) xor (A(101) and B(52)) xor (A(102) and B(51)) xor (A(103) and B(50)) xor (A(104) and B(49)) xor (A(105) and B(48)) xor (A(106) and B(47)) xor (A(107) and B(46)) xor (A(108) and B(45)) xor (A(109) and B(44)) xor (A(110) and B(43)) xor (A(111) and B(42)) xor (A(112) and B(41)) xor (A(113) and B(40)) xor (A(114) and B(39)) xor (A(115) and B(38)) xor (A(116) and B(37)) xor (A(117) and B(36)) xor (A(118) and B(35)) xor (A(119) and B(34)) xor (A(120) and B(33)) xor (A(121) and B(32)) xor (A(122) and B(31)) xor (A(123) and B(30)) xor (A(124) and B(29)) xor (A(125) and B(28)) xor (A(126) and B(28));
    C(27)  <= (A(0) and B(27)) xor (A(1) and B(26)) xor (A(2) and B(25)) xor (A(3) and B(24)) xor (A(4) and B(23)) xor (A(5) and B(23)) xor (A(6) and B(21)) xor (A(7) and B(20)) xor (A(8) and B(19)) xor (A(9) and B(18)) xor (A(10) and B(17)) xor (A(11) and B(16)) xor (A(12) and B(15)) xor (A(13) and B(14)) xor (A(14) and B(13)) xor (A(15) and B(12)) xor (A(16) and B(11)) xor (A(17) and B(10)) xor (A(18) and B(9)) xor (A(19) and B(8)) xor (A(20) and B(7)) xor (A(21) and B(6)) xor (A(23) and B(5)) xor (A(23) and B(4)) xor (A(24) and B(3)) xor (A(25) and B(2)) xor (A(26) and B(1)) xor (A(27) and B(0)) xor (A(20) and B(127)) xor (A(21) and B(126)) xor (A(23) and B(125)) xor (A(23) and B(124)) xor (A(24) and B(123)) xor (A(25) and B(122)) xor (A(26) and B(121)) xor (A(27) and B(120)) xor (A(28) and B(119)) xor (A(29) and B(118)) xor (A(30) and B(117)) xor (A(31) and B(116)) xor (A(32) and B(115)) xor (A(33) and B(114)) xor (A(34) and B(113)) xor (A(35) and B(112)) xor (A(36) and B(111)) xor (A(37) and B(110)) xor (A(38) and B(109)) xor (A(39) and B(108)) xor (A(40) and B(107)) xor (A(41) and B(106)) xor (A(42) and B(105)) xor (A(43) and B(104)) xor (A(44) and B(103)) xor (A(45) and B(102)) xor (A(46) and B(101)) xor (A(47) and B(100)) xor (A(48) and B(99)) xor (A(49) and B(98)) xor (A(50) and B(97)) xor (A(51) and B(96)) xor (A(52) and B(95)) xor (A(53) and B(94)) xor (A(54) and B(93)) xor (A(55) and B(92)) xor (A(56) and B(91)) xor (A(57) and B(90)) xor (A(58) and B(89)) xor (A(59) and B(88)) xor (A(60) and B(87)) xor (A(61) and B(86)) xor (A(62) and B(85)) xor (A(63) and B(84)) xor (A(64) and B(83)) xor (A(65) and B(82)) xor (A(66) and B(81)) xor (A(67) and B(80)) xor (A(68) and B(79)) xor (A(69) and B(78)) xor (A(70) and B(77)) xor (A(71) and B(76)) xor (A(72) and B(75)) xor (A(73) and B(74)) xor (A(74) and B(73)) xor (A(75) and B(72)) xor (A(76) and B(71)) xor (A(77) and B(70)) xor (A(78) and B(69)) xor (A(79) and B(68)) xor (A(80) and B(67)) xor (A(81) and B(66)) xor (A(82) and B(65)) xor (A(83) and B(64)) xor (A(84) and B(63)) xor (A(85) and B(62)) xor (A(86) and B(61)) xor (A(87) and B(60)) xor (A(88) and B(59)) xor (A(89) and B(58)) xor (A(90) and B(57)) xor (A(91) and B(56)) xor (A(92) and B(55)) xor (A(93) and B(54)) xor (A(94) and B(53)) xor (A(95) and B(52)) xor (A(96) and B(51)) xor (A(97) and B(50)) xor (A(98) and B(49)) xor (A(99) and B(48)) xor (A(100) and B(47)) xor (A(101) and B(46)) xor (A(102) and B(45)) xor (A(103) and B(44)) xor (A(104) and B(43)) xor (A(105) and B(42)) xor (A(106) and B(41)) xor (A(107) and B(40)) xor (A(108) and B(39)) xor (A(109) and B(38)) xor (A(110) and B(37)) xor (A(111) and B(36)) xor (A(112) and B(35)) xor (A(113) and B(34)) xor (A(114) and B(33)) xor (A(115) and B(32)) xor (A(116) and B(31)) xor (A(117) and B(30)) xor (A(118) and B(29)) xor (A(119) and B(28)) xor (A(120) and B(27)) xor (A(121) and B(26)) xor (A(122) and B(25)) xor (A(123) and B(24)) xor (A(124) and B(23)) xor (A(125) and B(23)) xor (A(126) and B(21)) xor (A(25) and B(127)) xor (A(26) and B(126)) xor (A(27) and B(125)) xor (A(28) and B(124)) xor (A(29) and B(123)) xor (A(30) and B(122)) xor (A(31) and B(121)) xor (A(32) and B(120)) xor (A(33) and B(119)) xor (A(34) and B(118)) xor (A(35) and B(117)) xor (A(36) and B(116)) xor (A(37) and B(115)) xor (A(38) and B(114)) xor (A(39) and B(113)) xor (A(40) and B(112)) xor (A(41) and B(111)) xor (A(42) and B(110)) xor (A(43) and B(109)) xor (A(44) and B(108)) xor (A(45) and B(107)) xor (A(46) and B(106)) xor (A(47) and B(105)) xor (A(48) and B(104)) xor (A(49) and B(103)) xor (A(50) and B(102)) xor (A(51) and B(101)) xor (A(52) and B(100)) xor (A(53) and B(99)) xor (A(54) and B(98)) xor (A(55) and B(97)) xor (A(56) and B(96)) xor (A(57) and B(95)) xor (A(58) and B(94)) xor (A(59) and B(93)) xor (A(60) and B(92)) xor (A(61) and B(91)) xor (A(62) and B(90)) xor (A(63) and B(89)) xor (A(64) and B(88)) xor (A(65) and B(87)) xor (A(66) and B(86)) xor (A(67) and B(85)) xor (A(68) and B(84)) xor (A(69) and B(83)) xor (A(70) and B(82)) xor (A(71) and B(81)) xor (A(72) and B(80)) xor (A(73) and B(79)) xor (A(74) and B(78)) xor (A(75) and B(77)) xor (A(76) and B(76)) xor (A(77) and B(75)) xor (A(78) and B(74)) xor (A(79) and B(73)) xor (A(80) and B(72)) xor (A(81) and B(71)) xor (A(82) and B(70)) xor (A(83) and B(69)) xor (A(84) and B(68)) xor (A(85) and B(67)) xor (A(86) and B(66)) xor (A(87) and B(65)) xor (A(88) and B(64)) xor (A(89) and B(63)) xor (A(90) and B(62)) xor (A(91) and B(61)) xor (A(92) and B(60)) xor (A(93) and B(59)) xor (A(94) and B(58)) xor (A(95) and B(57)) xor (A(96) and B(56)) xor (A(97) and B(55)) xor (A(98) and B(54)) xor (A(99) and B(53)) xor (A(100) and B(52)) xor (A(101) and B(51)) xor (A(102) and B(50)) xor (A(103) and B(49)) xor (A(104) and B(48)) xor (A(105) and B(47)) xor (A(106) and B(46)) xor (A(107) and B(45)) xor (A(108) and B(44)) xor (A(109) and B(43)) xor (A(110) and B(42)) xor (A(111) and B(41)) xor (A(112) and B(40)) xor (A(113) and B(39)) xor (A(114) and B(38)) xor (A(115) and B(37)) xor (A(116) and B(36)) xor (A(117) and B(35)) xor (A(118) and B(34)) xor (A(119) and B(33)) xor (A(120) and B(32)) xor (A(121) and B(31)) xor (A(122) and B(30)) xor (A(123) and B(29)) xor (A(124) and B(28)) xor (A(125) and B(27)) xor (A(126) and B(26)) xor (A(26) and B(127)) xor (A(27) and B(126)) xor (A(28) and B(125)) xor (A(29) and B(124)) xor (A(30) and B(123)) xor (A(31) and B(122)) xor (A(32) and B(121)) xor (A(33) and B(120)) xor (A(34) and B(119)) xor (A(35) and B(118)) xor (A(36) and B(117)) xor (A(37) and B(116)) xor (A(38) and B(115)) xor (A(39) and B(114)) xor (A(40) and B(113)) xor (A(41) and B(112)) xor (A(42) and B(111)) xor (A(43) and B(110)) xor (A(44) and B(109)) xor (A(45) and B(108)) xor (A(46) and B(107)) xor (A(47) and B(106)) xor (A(48) and B(105)) xor (A(49) and B(104)) xor (A(50) and B(103)) xor (A(51) and B(102)) xor (A(52) and B(101)) xor (A(53) and B(100)) xor (A(54) and B(99)) xor (A(55) and B(98)) xor (A(56) and B(97)) xor (A(57) and B(96)) xor (A(58) and B(95)) xor (A(59) and B(94)) xor (A(60) and B(93)) xor (A(61) and B(92)) xor (A(62) and B(91)) xor (A(63) and B(90)) xor (A(64) and B(89)) xor (A(65) and B(88)) xor (A(66) and B(87)) xor (A(67) and B(86)) xor (A(68) and B(85)) xor (A(69) and B(84)) xor (A(70) and B(83)) xor (A(71) and B(82)) xor (A(72) and B(81)) xor (A(73) and B(80)) xor (A(74) and B(79)) xor (A(75) and B(78)) xor (A(76) and B(77)) xor (A(77) and B(76)) xor (A(78) and B(75)) xor (A(79) and B(74)) xor (A(80) and B(73)) xor (A(81) and B(72)) xor (A(82) and B(71)) xor (A(83) and B(70)) xor (A(84) and B(69)) xor (A(85) and B(68)) xor (A(86) and B(67)) xor (A(87) and B(66)) xor (A(88) and B(65)) xor (A(89) and B(64)) xor (A(90) and B(63)) xor (A(91) and B(62)) xor (A(92) and B(61)) xor (A(93) and B(60)) xor (A(94) and B(59)) xor (A(95) and B(58)) xor (A(96) and B(57)) xor (A(97) and B(56)) xor (A(98) and B(55)) xor (A(99) and B(54)) xor (A(100) and B(53)) xor (A(101) and B(52)) xor (A(102) and B(51)) xor (A(103) and B(50)) xor (A(104) and B(49)) xor (A(105) and B(48)) xor (A(106) and B(47)) xor (A(107) and B(46)) xor (A(108) and B(45)) xor (A(109) and B(44)) xor (A(110) and B(43)) xor (A(111) and B(42)) xor (A(112) and B(41)) xor (A(113) and B(40)) xor (A(114) and B(39)) xor (A(115) and B(38)) xor (A(116) and B(37)) xor (A(117) and B(36)) xor (A(118) and B(35)) xor (A(119) and B(34)) xor (A(120) and B(33)) xor (A(121) and B(32)) xor (A(122) and B(31)) xor (A(123) and B(30)) xor (A(124) and B(29)) xor (A(125) and B(28)) xor (A(126) and B(27)) xor (A(27) and B(127)) xor (A(28) and B(126)) xor (A(29) and B(125)) xor (A(30) and B(124)) xor (A(31) and B(123)) xor (A(32) and B(122)) xor (A(33) and B(121)) xor (A(34) and B(120)) xor (A(35) and B(119)) xor (A(36) and B(118)) xor (A(37) and B(117)) xor (A(38) and B(116)) xor (A(39) and B(115)) xor (A(40) and B(114)) xor (A(41) and B(113)) xor (A(42) and B(112)) xor (A(43) and B(111)) xor (A(44) and B(110)) xor (A(45) and B(109)) xor (A(46) and B(108)) xor (A(47) and B(107)) xor (A(48) and B(106)) xor (A(49) and B(105)) xor (A(50) and B(104)) xor (A(51) and B(103)) xor (A(52) and B(102)) xor (A(53) and B(101)) xor (A(54) and B(100)) xor (A(55) and B(99)) xor (A(56) and B(98)) xor (A(57) and B(97)) xor (A(58) and B(96)) xor (A(59) and B(95)) xor (A(60) and B(94)) xor (A(61) and B(93)) xor (A(62) and B(92)) xor (A(63) and B(91)) xor (A(64) and B(90)) xor (A(65) and B(89)) xor (A(66) and B(88)) xor (A(67) and B(87)) xor (A(68) and B(86)) xor (A(69) and B(85)) xor (A(70) and B(84)) xor (A(71) and B(83)) xor (A(72) and B(82)) xor (A(73) and B(81)) xor (A(74) and B(80)) xor (A(75) and B(79)) xor (A(76) and B(78)) xor (A(77) and B(77)) xor (A(78) and B(76)) xor (A(79) and B(75)) xor (A(80) and B(74)) xor (A(81) and B(73)) xor (A(82) and B(72)) xor (A(83) and B(71)) xor (A(84) and B(70)) xor (A(85) and B(69)) xor (A(86) and B(68)) xor (A(87) and B(67)) xor (A(88) and B(66)) xor (A(89) and B(65)) xor (A(90) and B(64)) xor (A(91) and B(63)) xor (A(92) and B(62)) xor (A(93) and B(61)) xor (A(94) and B(60)) xor (A(95) and B(59)) xor (A(96) and B(58)) xor (A(97) and B(57)) xor (A(98) and B(56)) xor (A(99) and B(55)) xor (A(100) and B(54)) xor (A(101) and B(53)) xor (A(102) and B(52)) xor (A(103) and B(51)) xor (A(104) and B(50)) xor (A(105) and B(49)) xor (A(106) and B(48)) xor (A(107) and B(47)) xor (A(108) and B(46)) xor (A(109) and B(45)) xor (A(110) and B(44)) xor (A(111) and B(43)) xor (A(112) and B(42)) xor (A(113) and B(41)) xor (A(114) and B(40)) xor (A(115) and B(39)) xor (A(116) and B(38)) xor (A(117) and B(37)) xor (A(118) and B(36)) xor (A(119) and B(35)) xor (A(120) and B(34)) xor (A(121) and B(33)) xor (A(122) and B(32)) xor (A(123) and B(31)) xor (A(124) and B(30)) xor (A(125) and B(29)) xor (A(126) and B(29));
    C(28)  <= (A(0) and B(28)) xor (A(1) and B(27)) xor (A(2) and B(26)) xor (A(3) and B(25)) xor (A(4) and B(24)) xor (A(5) and B(23)) xor (A(6) and B(23)) xor (A(7) and B(21)) xor (A(8) and B(20)) xor (A(9) and B(19)) xor (A(10) and B(18)) xor (A(11) and B(17)) xor (A(12) and B(16)) xor (A(13) and B(15)) xor (A(14) and B(14)) xor (A(15) and B(13)) xor (A(16) and B(12)) xor (A(17) and B(11)) xor (A(18) and B(10)) xor (A(19) and B(9)) xor (A(20) and B(8)) xor (A(21) and B(7)) xor (A(23) and B(6)) xor (A(23) and B(5)) xor (A(24) and B(4)) xor (A(25) and B(3)) xor (A(26) and B(2)) xor (A(27) and B(1)) xor (A(28) and B(0)) xor (A(21) and B(127)) xor (A(23) and B(126)) xor (A(23) and B(125)) xor (A(24) and B(124)) xor (A(25) and B(123)) xor (A(26) and B(122)) xor (A(27) and B(121)) xor (A(28) and B(120)) xor (A(29) and B(119)) xor (A(30) and B(118)) xor (A(31) and B(117)) xor (A(32) and B(116)) xor (A(33) and B(115)) xor (A(34) and B(114)) xor (A(35) and B(113)) xor (A(36) and B(112)) xor (A(37) and B(111)) xor (A(38) and B(110)) xor (A(39) and B(109)) xor (A(40) and B(108)) xor (A(41) and B(107)) xor (A(42) and B(106)) xor (A(43) and B(105)) xor (A(44) and B(104)) xor (A(45) and B(103)) xor (A(46) and B(102)) xor (A(47) and B(101)) xor (A(48) and B(100)) xor (A(49) and B(99)) xor (A(50) and B(98)) xor (A(51) and B(97)) xor (A(52) and B(96)) xor (A(53) and B(95)) xor (A(54) and B(94)) xor (A(55) and B(93)) xor (A(56) and B(92)) xor (A(57) and B(91)) xor (A(58) and B(90)) xor (A(59) and B(89)) xor (A(60) and B(88)) xor (A(61) and B(87)) xor (A(62) and B(86)) xor (A(63) and B(85)) xor (A(64) and B(84)) xor (A(65) and B(83)) xor (A(66) and B(82)) xor (A(67) and B(81)) xor (A(68) and B(80)) xor (A(69) and B(79)) xor (A(70) and B(78)) xor (A(71) and B(77)) xor (A(72) and B(76)) xor (A(73) and B(75)) xor (A(74) and B(74)) xor (A(75) and B(73)) xor (A(76) and B(72)) xor (A(77) and B(71)) xor (A(78) and B(70)) xor (A(79) and B(69)) xor (A(80) and B(68)) xor (A(81) and B(67)) xor (A(82) and B(66)) xor (A(83) and B(65)) xor (A(84) and B(64)) xor (A(85) and B(63)) xor (A(86) and B(62)) xor (A(87) and B(61)) xor (A(88) and B(60)) xor (A(89) and B(59)) xor (A(90) and B(58)) xor (A(91) and B(57)) xor (A(92) and B(56)) xor (A(93) and B(55)) xor (A(94) and B(54)) xor (A(95) and B(53)) xor (A(96) and B(52)) xor (A(97) and B(51)) xor (A(98) and B(50)) xor (A(99) and B(49)) xor (A(100) and B(48)) xor (A(101) and B(47)) xor (A(102) and B(46)) xor (A(103) and B(45)) xor (A(104) and B(44)) xor (A(105) and B(43)) xor (A(106) and B(42)) xor (A(107) and B(41)) xor (A(108) and B(40)) xor (A(109) and B(39)) xor (A(110) and B(38)) xor (A(111) and B(37)) xor (A(112) and B(36)) xor (A(113) and B(35)) xor (A(114) and B(34)) xor (A(115) and B(33)) xor (A(116) and B(32)) xor (A(117) and B(31)) xor (A(118) and B(30)) xor (A(119) and B(29)) xor (A(120) and B(28)) xor (A(121) and B(27)) xor (A(122) and B(26)) xor (A(123) and B(25)) xor (A(124) and B(24)) xor (A(125) and B(23)) xor (A(126) and B(23)) xor (A(26) and B(127)) xor (A(27) and B(126)) xor (A(28) and B(125)) xor (A(29) and B(124)) xor (A(30) and B(123)) xor (A(31) and B(122)) xor (A(32) and B(121)) xor (A(33) and B(120)) xor (A(34) and B(119)) xor (A(35) and B(118)) xor (A(36) and B(117)) xor (A(37) and B(116)) xor (A(38) and B(115)) xor (A(39) and B(114)) xor (A(40) and B(113)) xor (A(41) and B(112)) xor (A(42) and B(111)) xor (A(43) and B(110)) xor (A(44) and B(109)) xor (A(45) and B(108)) xor (A(46) and B(107)) xor (A(47) and B(106)) xor (A(48) and B(105)) xor (A(49) and B(104)) xor (A(50) and B(103)) xor (A(51) and B(102)) xor (A(52) and B(101)) xor (A(53) and B(100)) xor (A(54) and B(99)) xor (A(55) and B(98)) xor (A(56) and B(97)) xor (A(57) and B(96)) xor (A(58) and B(95)) xor (A(59) and B(94)) xor (A(60) and B(93)) xor (A(61) and B(92)) xor (A(62) and B(91)) xor (A(63) and B(90)) xor (A(64) and B(89)) xor (A(65) and B(88)) xor (A(66) and B(87)) xor (A(67) and B(86)) xor (A(68) and B(85)) xor (A(69) and B(84)) xor (A(70) and B(83)) xor (A(71) and B(82)) xor (A(72) and B(81)) xor (A(73) and B(80)) xor (A(74) and B(79)) xor (A(75) and B(78)) xor (A(76) and B(77)) xor (A(77) and B(76)) xor (A(78) and B(75)) xor (A(79) and B(74)) xor (A(80) and B(73)) xor (A(81) and B(72)) xor (A(82) and B(71)) xor (A(83) and B(70)) xor (A(84) and B(69)) xor (A(85) and B(68)) xor (A(86) and B(67)) xor (A(87) and B(66)) xor (A(88) and B(65)) xor (A(89) and B(64)) xor (A(90) and B(63)) xor (A(91) and B(62)) xor (A(92) and B(61)) xor (A(93) and B(60)) xor (A(94) and B(59)) xor (A(95) and B(58)) xor (A(96) and B(57)) xor (A(97) and B(56)) xor (A(98) and B(55)) xor (A(99) and B(54)) xor (A(100) and B(53)) xor (A(101) and B(52)) xor (A(102) and B(51)) xor (A(103) and B(50)) xor (A(104) and B(49)) xor (A(105) and B(48)) xor (A(106) and B(47)) xor (A(107) and B(46)) xor (A(108) and B(45)) xor (A(109) and B(44)) xor (A(110) and B(43)) xor (A(111) and B(42)) xor (A(112) and B(41)) xor (A(113) and B(40)) xor (A(114) and B(39)) xor (A(115) and B(38)) xor (A(116) and B(37)) xor (A(117) and B(36)) xor (A(118) and B(35)) xor (A(119) and B(34)) xor (A(120) and B(33)) xor (A(121) and B(32)) xor (A(122) and B(31)) xor (A(123) and B(30)) xor (A(124) and B(29)) xor (A(125) and B(28)) xor (A(126) and B(27)) xor (A(27) and B(127)) xor (A(28) and B(126)) xor (A(29) and B(125)) xor (A(30) and B(124)) xor (A(31) and B(123)) xor (A(32) and B(122)) xor (A(33) and B(121)) xor (A(34) and B(120)) xor (A(35) and B(119)) xor (A(36) and B(118)) xor (A(37) and B(117)) xor (A(38) and B(116)) xor (A(39) and B(115)) xor (A(40) and B(114)) xor (A(41) and B(113)) xor (A(42) and B(112)) xor (A(43) and B(111)) xor (A(44) and B(110)) xor (A(45) and B(109)) xor (A(46) and B(108)) xor (A(47) and B(107)) xor (A(48) and B(106)) xor (A(49) and B(105)) xor (A(50) and B(104)) xor (A(51) and B(103)) xor (A(52) and B(102)) xor (A(53) and B(101)) xor (A(54) and B(100)) xor (A(55) and B(99)) xor (A(56) and B(98)) xor (A(57) and B(97)) xor (A(58) and B(96)) xor (A(59) and B(95)) xor (A(60) and B(94)) xor (A(61) and B(93)) xor (A(62) and B(92)) xor (A(63) and B(91)) xor (A(64) and B(90)) xor (A(65) and B(89)) xor (A(66) and B(88)) xor (A(67) and B(87)) xor (A(68) and B(86)) xor (A(69) and B(85)) xor (A(70) and B(84)) xor (A(71) and B(83)) xor (A(72) and B(82)) xor (A(73) and B(81)) xor (A(74) and B(80)) xor (A(75) and B(79)) xor (A(76) and B(78)) xor (A(77) and B(77)) xor (A(78) and B(76)) xor (A(79) and B(75)) xor (A(80) and B(74)) xor (A(81) and B(73)) xor (A(82) and B(72)) xor (A(83) and B(71)) xor (A(84) and B(70)) xor (A(85) and B(69)) xor (A(86) and B(68)) xor (A(87) and B(67)) xor (A(88) and B(66)) xor (A(89) and B(65)) xor (A(90) and B(64)) xor (A(91) and B(63)) xor (A(92) and B(62)) xor (A(93) and B(61)) xor (A(94) and B(60)) xor (A(95) and B(59)) xor (A(96) and B(58)) xor (A(97) and B(57)) xor (A(98) and B(56)) xor (A(99) and B(55)) xor (A(100) and B(54)) xor (A(101) and B(53)) xor (A(102) and B(52)) xor (A(103) and B(51)) xor (A(104) and B(50)) xor (A(105) and B(49)) xor (A(106) and B(48)) xor (A(107) and B(47)) xor (A(108) and B(46)) xor (A(109) and B(45)) xor (A(110) and B(44)) xor (A(111) and B(43)) xor (A(112) and B(42)) xor (A(113) and B(41)) xor (A(114) and B(40)) xor (A(115) and B(39)) xor (A(116) and B(38)) xor (A(117) and B(37)) xor (A(118) and B(36)) xor (A(119) and B(35)) xor (A(120) and B(34)) xor (A(121) and B(33)) xor (A(122) and B(32)) xor (A(123) and B(31)) xor (A(124) and B(30)) xor (A(125) and B(29)) xor (A(126) and B(28)) xor (A(28) and B(127)) xor (A(29) and B(126)) xor (A(30) and B(125)) xor (A(31) and B(124)) xor (A(32) and B(123)) xor (A(33) and B(122)) xor (A(34) and B(121)) xor (A(35) and B(120)) xor (A(36) and B(119)) xor (A(37) and B(118)) xor (A(38) and B(117)) xor (A(39) and B(116)) xor (A(40) and B(115)) xor (A(41) and B(114)) xor (A(42) and B(113)) xor (A(43) and B(112)) xor (A(44) and B(111)) xor (A(45) and B(110)) xor (A(46) and B(109)) xor (A(47) and B(108)) xor (A(48) and B(107)) xor (A(49) and B(106)) xor (A(50) and B(105)) xor (A(51) and B(104)) xor (A(52) and B(103)) xor (A(53) and B(102)) xor (A(54) and B(101)) xor (A(55) and B(100)) xor (A(56) and B(99)) xor (A(57) and B(98)) xor (A(58) and B(97)) xor (A(59) and B(96)) xor (A(60) and B(95)) xor (A(61) and B(94)) xor (A(62) and B(93)) xor (A(63) and B(92)) xor (A(64) and B(91)) xor (A(65) and B(90)) xor (A(66) and B(89)) xor (A(67) and B(88)) xor (A(68) and B(87)) xor (A(69) and B(86)) xor (A(70) and B(85)) xor (A(71) and B(84)) xor (A(72) and B(83)) xor (A(73) and B(82)) xor (A(74) and B(81)) xor (A(75) and B(80)) xor (A(76) and B(79)) xor (A(77) and B(78)) xor (A(78) and B(77)) xor (A(79) and B(76)) xor (A(80) and B(75)) xor (A(81) and B(74)) xor (A(82) and B(73)) xor (A(83) and B(72)) xor (A(84) and B(71)) xor (A(85) and B(70)) xor (A(86) and B(69)) xor (A(87) and B(68)) xor (A(88) and B(67)) xor (A(89) and B(66)) xor (A(90) and B(65)) xor (A(91) and B(64)) xor (A(92) and B(63)) xor (A(93) and B(62)) xor (A(94) and B(61)) xor (A(95) and B(60)) xor (A(96) and B(59)) xor (A(97) and B(58)) xor (A(98) and B(57)) xor (A(99) and B(56)) xor (A(100) and B(55)) xor (A(101) and B(54)) xor (A(102) and B(53)) xor (A(103) and B(52)) xor (A(104) and B(51)) xor (A(105) and B(50)) xor (A(106) and B(49)) xor (A(107) and B(48)) xor (A(108) and B(47)) xor (A(109) and B(46)) xor (A(110) and B(45)) xor (A(111) and B(44)) xor (A(112) and B(43)) xor (A(113) and B(42)) xor (A(114) and B(41)) xor (A(115) and B(40)) xor (A(116) and B(39)) xor (A(117) and B(38)) xor (A(118) and B(37)) xor (A(119) and B(36)) xor (A(120) and B(35)) xor (A(121) and B(34)) xor (A(122) and B(33)) xor (A(123) and B(32)) xor (A(124) and B(31)) xor (A(125) and B(30)) xor (A(126) and B(30));
    C(29)  <= (A(0) and B(29)) xor (A(1) and B(28)) xor (A(2) and B(27)) xor (A(3) and B(26)) xor (A(4) and B(25)) xor (A(5) and B(24)) xor (A(6) and B(23)) xor (A(7) and B(23)) xor (A(8) and B(21)) xor (A(9) and B(20)) xor (A(10) and B(19)) xor (A(11) and B(18)) xor (A(12) and B(17)) xor (A(13) and B(16)) xor (A(14) and B(15)) xor (A(15) and B(14)) xor (A(16) and B(13)) xor (A(17) and B(12)) xor (A(18) and B(11)) xor (A(19) and B(10)) xor (A(20) and B(9)) xor (A(21) and B(8)) xor (A(23) and B(7)) xor (A(23) and B(6)) xor (A(24) and B(5)) xor (A(25) and B(4)) xor (A(26) and B(3)) xor (A(27) and B(2)) xor (A(28) and B(1)) xor (A(29) and B(0)) xor (A(23) and B(127)) xor (A(23) and B(126)) xor (A(24) and B(125)) xor (A(25) and B(124)) xor (A(26) and B(123)) xor (A(27) and B(122)) xor (A(28) and B(121)) xor (A(29) and B(120)) xor (A(30) and B(119)) xor (A(31) and B(118)) xor (A(32) and B(117)) xor (A(33) and B(116)) xor (A(34) and B(115)) xor (A(35) and B(114)) xor (A(36) and B(113)) xor (A(37) and B(112)) xor (A(38) and B(111)) xor (A(39) and B(110)) xor (A(40) and B(109)) xor (A(41) and B(108)) xor (A(42) and B(107)) xor (A(43) and B(106)) xor (A(44) and B(105)) xor (A(45) and B(104)) xor (A(46) and B(103)) xor (A(47) and B(102)) xor (A(48) and B(101)) xor (A(49) and B(100)) xor (A(50) and B(99)) xor (A(51) and B(98)) xor (A(52) and B(97)) xor (A(53) and B(96)) xor (A(54) and B(95)) xor (A(55) and B(94)) xor (A(56) and B(93)) xor (A(57) and B(92)) xor (A(58) and B(91)) xor (A(59) and B(90)) xor (A(60) and B(89)) xor (A(61) and B(88)) xor (A(62) and B(87)) xor (A(63) and B(86)) xor (A(64) and B(85)) xor (A(65) and B(84)) xor (A(66) and B(83)) xor (A(67) and B(82)) xor (A(68) and B(81)) xor (A(69) and B(80)) xor (A(70) and B(79)) xor (A(71) and B(78)) xor (A(72) and B(77)) xor (A(73) and B(76)) xor (A(74) and B(75)) xor (A(75) and B(74)) xor (A(76) and B(73)) xor (A(77) and B(72)) xor (A(78) and B(71)) xor (A(79) and B(70)) xor (A(80) and B(69)) xor (A(81) and B(68)) xor (A(82) and B(67)) xor (A(83) and B(66)) xor (A(84) and B(65)) xor (A(85) and B(64)) xor (A(86) and B(63)) xor (A(87) and B(62)) xor (A(88) and B(61)) xor (A(89) and B(60)) xor (A(90) and B(59)) xor (A(91) and B(58)) xor (A(92) and B(57)) xor (A(93) and B(56)) xor (A(94) and B(55)) xor (A(95) and B(54)) xor (A(96) and B(53)) xor (A(97) and B(52)) xor (A(98) and B(51)) xor (A(99) and B(50)) xor (A(100) and B(49)) xor (A(101) and B(48)) xor (A(102) and B(47)) xor (A(103) and B(46)) xor (A(104) and B(45)) xor (A(105) and B(44)) xor (A(106) and B(43)) xor (A(107) and B(42)) xor (A(108) and B(41)) xor (A(109) and B(40)) xor (A(110) and B(39)) xor (A(111) and B(38)) xor (A(112) and B(37)) xor (A(113) and B(36)) xor (A(114) and B(35)) xor (A(115) and B(34)) xor (A(116) and B(33)) xor (A(117) and B(32)) xor (A(118) and B(31)) xor (A(119) and B(30)) xor (A(120) and B(29)) xor (A(121) and B(28)) xor (A(122) and B(27)) xor (A(123) and B(26)) xor (A(124) and B(25)) xor (A(125) and B(24)) xor (A(126) and B(23)) xor (A(27) and B(127)) xor (A(28) and B(126)) xor (A(29) and B(125)) xor (A(30) and B(124)) xor (A(31) and B(123)) xor (A(32) and B(122)) xor (A(33) and B(121)) xor (A(34) and B(120)) xor (A(35) and B(119)) xor (A(36) and B(118)) xor (A(37) and B(117)) xor (A(38) and B(116)) xor (A(39) and B(115)) xor (A(40) and B(114)) xor (A(41) and B(113)) xor (A(42) and B(112)) xor (A(43) and B(111)) xor (A(44) and B(110)) xor (A(45) and B(109)) xor (A(46) and B(108)) xor (A(47) and B(107)) xor (A(48) and B(106)) xor (A(49) and B(105)) xor (A(50) and B(104)) xor (A(51) and B(103)) xor (A(52) and B(102)) xor (A(53) and B(101)) xor (A(54) and B(100)) xor (A(55) and B(99)) xor (A(56) and B(98)) xor (A(57) and B(97)) xor (A(58) and B(96)) xor (A(59) and B(95)) xor (A(60) and B(94)) xor (A(61) and B(93)) xor (A(62) and B(92)) xor (A(63) and B(91)) xor (A(64) and B(90)) xor (A(65) and B(89)) xor (A(66) and B(88)) xor (A(67) and B(87)) xor (A(68) and B(86)) xor (A(69) and B(85)) xor (A(70) and B(84)) xor (A(71) and B(83)) xor (A(72) and B(82)) xor (A(73) and B(81)) xor (A(74) and B(80)) xor (A(75) and B(79)) xor (A(76) and B(78)) xor (A(77) and B(77)) xor (A(78) and B(76)) xor (A(79) and B(75)) xor (A(80) and B(74)) xor (A(81) and B(73)) xor (A(82) and B(72)) xor (A(83) and B(71)) xor (A(84) and B(70)) xor (A(85) and B(69)) xor (A(86) and B(68)) xor (A(87) and B(67)) xor (A(88) and B(66)) xor (A(89) and B(65)) xor (A(90) and B(64)) xor (A(91) and B(63)) xor (A(92) and B(62)) xor (A(93) and B(61)) xor (A(94) and B(60)) xor (A(95) and B(59)) xor (A(96) and B(58)) xor (A(97) and B(57)) xor (A(98) and B(56)) xor (A(99) and B(55)) xor (A(100) and B(54)) xor (A(101) and B(53)) xor (A(102) and B(52)) xor (A(103) and B(51)) xor (A(104) and B(50)) xor (A(105) and B(49)) xor (A(106) and B(48)) xor (A(107) and B(47)) xor (A(108) and B(46)) xor (A(109) and B(45)) xor (A(110) and B(44)) xor (A(111) and B(43)) xor (A(112) and B(42)) xor (A(113) and B(41)) xor (A(114) and B(40)) xor (A(115) and B(39)) xor (A(116) and B(38)) xor (A(117) and B(37)) xor (A(118) and B(36)) xor (A(119) and B(35)) xor (A(120) and B(34)) xor (A(121) and B(33)) xor (A(122) and B(32)) xor (A(123) and B(31)) xor (A(124) and B(30)) xor (A(125) and B(29)) xor (A(126) and B(28)) xor (A(28) and B(127)) xor (A(29) and B(126)) xor (A(30) and B(125)) xor (A(31) and B(124)) xor (A(32) and B(123)) xor (A(33) and B(122)) xor (A(34) and B(121)) xor (A(35) and B(120)) xor (A(36) and B(119)) xor (A(37) and B(118)) xor (A(38) and B(117)) xor (A(39) and B(116)) xor (A(40) and B(115)) xor (A(41) and B(114)) xor (A(42) and B(113)) xor (A(43) and B(112)) xor (A(44) and B(111)) xor (A(45) and B(110)) xor (A(46) and B(109)) xor (A(47) and B(108)) xor (A(48) and B(107)) xor (A(49) and B(106)) xor (A(50) and B(105)) xor (A(51) and B(104)) xor (A(52) and B(103)) xor (A(53) and B(102)) xor (A(54) and B(101)) xor (A(55) and B(100)) xor (A(56) and B(99)) xor (A(57) and B(98)) xor (A(58) and B(97)) xor (A(59) and B(96)) xor (A(60) and B(95)) xor (A(61) and B(94)) xor (A(62) and B(93)) xor (A(63) and B(92)) xor (A(64) and B(91)) xor (A(65) and B(90)) xor (A(66) and B(89)) xor (A(67) and B(88)) xor (A(68) and B(87)) xor (A(69) and B(86)) xor (A(70) and B(85)) xor (A(71) and B(84)) xor (A(72) and B(83)) xor (A(73) and B(82)) xor (A(74) and B(81)) xor (A(75) and B(80)) xor (A(76) and B(79)) xor (A(77) and B(78)) xor (A(78) and B(77)) xor (A(79) and B(76)) xor (A(80) and B(75)) xor (A(81) and B(74)) xor (A(82) and B(73)) xor (A(83) and B(72)) xor (A(84) and B(71)) xor (A(85) and B(70)) xor (A(86) and B(69)) xor (A(87) and B(68)) xor (A(88) and B(67)) xor (A(89) and B(66)) xor (A(90) and B(65)) xor (A(91) and B(64)) xor (A(92) and B(63)) xor (A(93) and B(62)) xor (A(94) and B(61)) xor (A(95) and B(60)) xor (A(96) and B(59)) xor (A(97) and B(58)) xor (A(98) and B(57)) xor (A(99) and B(56)) xor (A(100) and B(55)) xor (A(101) and B(54)) xor (A(102) and B(53)) xor (A(103) and B(52)) xor (A(104) and B(51)) xor (A(105) and B(50)) xor (A(106) and B(49)) xor (A(107) and B(48)) xor (A(108) and B(47)) xor (A(109) and B(46)) xor (A(110) and B(45)) xor (A(111) and B(44)) xor (A(112) and B(43)) xor (A(113) and B(42)) xor (A(114) and B(41)) xor (A(115) and B(40)) xor (A(116) and B(39)) xor (A(117) and B(38)) xor (A(118) and B(37)) xor (A(119) and B(36)) xor (A(120) and B(35)) xor (A(121) and B(34)) xor (A(122) and B(33)) xor (A(123) and B(32)) xor (A(124) and B(31)) xor (A(125) and B(30)) xor (A(126) and B(29)) xor (A(29) and B(127)) xor (A(30) and B(126)) xor (A(31) and B(125)) xor (A(32) and B(124)) xor (A(33) and B(123)) xor (A(34) and B(122)) xor (A(35) and B(121)) xor (A(36) and B(120)) xor (A(37) and B(119)) xor (A(38) and B(118)) xor (A(39) and B(117)) xor (A(40) and B(116)) xor (A(41) and B(115)) xor (A(42) and B(114)) xor (A(43) and B(113)) xor (A(44) and B(112)) xor (A(45) and B(111)) xor (A(46) and B(110)) xor (A(47) and B(109)) xor (A(48) and B(108)) xor (A(49) and B(107)) xor (A(50) and B(106)) xor (A(51) and B(105)) xor (A(52) and B(104)) xor (A(53) and B(103)) xor (A(54) and B(102)) xor (A(55) and B(101)) xor (A(56) and B(100)) xor (A(57) and B(99)) xor (A(58) and B(98)) xor (A(59) and B(97)) xor (A(60) and B(96)) xor (A(61) and B(95)) xor (A(62) and B(94)) xor (A(63) and B(93)) xor (A(64) and B(92)) xor (A(65) and B(91)) xor (A(66) and B(90)) xor (A(67) and B(89)) xor (A(68) and B(88)) xor (A(69) and B(87)) xor (A(70) and B(86)) xor (A(71) and B(85)) xor (A(72) and B(84)) xor (A(73) and B(83)) xor (A(74) and B(82)) xor (A(75) and B(81)) xor (A(76) and B(80)) xor (A(77) and B(79)) xor (A(78) and B(78)) xor (A(79) and B(77)) xor (A(80) and B(76)) xor (A(81) and B(75)) xor (A(82) and B(74)) xor (A(83) and B(73)) xor (A(84) and B(72)) xor (A(85) and B(71)) xor (A(86) and B(70)) xor (A(87) and B(69)) xor (A(88) and B(68)) xor (A(89) and B(67)) xor (A(90) and B(66)) xor (A(91) and B(65)) xor (A(92) and B(64)) xor (A(93) and B(63)) xor (A(94) and B(62)) xor (A(95) and B(61)) xor (A(96) and B(60)) xor (A(97) and B(59)) xor (A(98) and B(58)) xor (A(99) and B(57)) xor (A(100) and B(56)) xor (A(101) and B(55)) xor (A(102) and B(54)) xor (A(103) and B(53)) xor (A(104) and B(52)) xor (A(105) and B(51)) xor (A(106) and B(50)) xor (A(107) and B(49)) xor (A(108) and B(48)) xor (A(109) and B(47)) xor (A(110) and B(46)) xor (A(111) and B(45)) xor (A(112) and B(44)) xor (A(113) and B(43)) xor (A(114) and B(42)) xor (A(115) and B(41)) xor (A(116) and B(40)) xor (A(117) and B(39)) xor (A(118) and B(38)) xor (A(119) and B(37)) xor (A(120) and B(36)) xor (A(121) and B(35)) xor (A(122) and B(34)) xor (A(123) and B(33)) xor (A(124) and B(32)) xor (A(125) and B(31)) xor (A(126) and B(31));
    C(30)  <= (A(0) and B(30)) xor (A(1) and B(29)) xor (A(2) and B(28)) xor (A(3) and B(27)) xor (A(4) and B(26)) xor (A(5) and B(25)) xor (A(6) and B(24)) xor (A(7) and B(23)) xor (A(8) and B(23)) xor (A(9) and B(21)) xor (A(10) and B(20)) xor (A(11) and B(19)) xor (A(12) and B(18)) xor (A(13) and B(17)) xor (A(14) and B(16)) xor (A(15) and B(15)) xor (A(16) and B(14)) xor (A(17) and B(13)) xor (A(18) and B(12)) xor (A(19) and B(11)) xor (A(20) and B(10)) xor (A(21) and B(9)) xor (A(23) and B(8)) xor (A(23) and B(7)) xor (A(24) and B(6)) xor (A(25) and B(5)) xor (A(26) and B(4)) xor (A(27) and B(3)) xor (A(28) and B(2)) xor (A(29) and B(1)) xor (A(30) and B(0)) xor (A(23) and B(127)) xor (A(24) and B(126)) xor (A(25) and B(125)) xor (A(26) and B(124)) xor (A(27) and B(123)) xor (A(28) and B(122)) xor (A(29) and B(121)) xor (A(30) and B(120)) xor (A(31) and B(119)) xor (A(32) and B(118)) xor (A(33) and B(117)) xor (A(34) and B(116)) xor (A(35) and B(115)) xor (A(36) and B(114)) xor (A(37) and B(113)) xor (A(38) and B(112)) xor (A(39) and B(111)) xor (A(40) and B(110)) xor (A(41) and B(109)) xor (A(42) and B(108)) xor (A(43) and B(107)) xor (A(44) and B(106)) xor (A(45) and B(105)) xor (A(46) and B(104)) xor (A(47) and B(103)) xor (A(48) and B(102)) xor (A(49) and B(101)) xor (A(50) and B(100)) xor (A(51) and B(99)) xor (A(52) and B(98)) xor (A(53) and B(97)) xor (A(54) and B(96)) xor (A(55) and B(95)) xor (A(56) and B(94)) xor (A(57) and B(93)) xor (A(58) and B(92)) xor (A(59) and B(91)) xor (A(60) and B(90)) xor (A(61) and B(89)) xor (A(62) and B(88)) xor (A(63) and B(87)) xor (A(64) and B(86)) xor (A(65) and B(85)) xor (A(66) and B(84)) xor (A(67) and B(83)) xor (A(68) and B(82)) xor (A(69) and B(81)) xor (A(70) and B(80)) xor (A(71) and B(79)) xor (A(72) and B(78)) xor (A(73) and B(77)) xor (A(74) and B(76)) xor (A(75) and B(75)) xor (A(76) and B(74)) xor (A(77) and B(73)) xor (A(78) and B(72)) xor (A(79) and B(71)) xor (A(80) and B(70)) xor (A(81) and B(69)) xor (A(82) and B(68)) xor (A(83) and B(67)) xor (A(84) and B(66)) xor (A(85) and B(65)) xor (A(86) and B(64)) xor (A(87) and B(63)) xor (A(88) and B(62)) xor (A(89) and B(61)) xor (A(90) and B(60)) xor (A(91) and B(59)) xor (A(92) and B(58)) xor (A(93) and B(57)) xor (A(94) and B(56)) xor (A(95) and B(55)) xor (A(96) and B(54)) xor (A(97) and B(53)) xor (A(98) and B(52)) xor (A(99) and B(51)) xor (A(100) and B(50)) xor (A(101) and B(49)) xor (A(102) and B(48)) xor (A(103) and B(47)) xor (A(104) and B(46)) xor (A(105) and B(45)) xor (A(106) and B(44)) xor (A(107) and B(43)) xor (A(108) and B(42)) xor (A(109) and B(41)) xor (A(110) and B(40)) xor (A(111) and B(39)) xor (A(112) and B(38)) xor (A(113) and B(37)) xor (A(114) and B(36)) xor (A(115) and B(35)) xor (A(116) and B(34)) xor (A(117) and B(33)) xor (A(118) and B(32)) xor (A(119) and B(31)) xor (A(120) and B(30)) xor (A(121) and B(29)) xor (A(122) and B(28)) xor (A(123) and B(27)) xor (A(124) and B(26)) xor (A(125) and B(25)) xor (A(126) and B(24)) xor (A(28) and B(127)) xor (A(29) and B(126)) xor (A(30) and B(125)) xor (A(31) and B(124)) xor (A(32) and B(123)) xor (A(33) and B(122)) xor (A(34) and B(121)) xor (A(35) and B(120)) xor (A(36) and B(119)) xor (A(37) and B(118)) xor (A(38) and B(117)) xor (A(39) and B(116)) xor (A(40) and B(115)) xor (A(41) and B(114)) xor (A(42) and B(113)) xor (A(43) and B(112)) xor (A(44) and B(111)) xor (A(45) and B(110)) xor (A(46) and B(109)) xor (A(47) and B(108)) xor (A(48) and B(107)) xor (A(49) and B(106)) xor (A(50) and B(105)) xor (A(51) and B(104)) xor (A(52) and B(103)) xor (A(53) and B(102)) xor (A(54) and B(101)) xor (A(55) and B(100)) xor (A(56) and B(99)) xor (A(57) and B(98)) xor (A(58) and B(97)) xor (A(59) and B(96)) xor (A(60) and B(95)) xor (A(61) and B(94)) xor (A(62) and B(93)) xor (A(63) and B(92)) xor (A(64) and B(91)) xor (A(65) and B(90)) xor (A(66) and B(89)) xor (A(67) and B(88)) xor (A(68) and B(87)) xor (A(69) and B(86)) xor (A(70) and B(85)) xor (A(71) and B(84)) xor (A(72) and B(83)) xor (A(73) and B(82)) xor (A(74) and B(81)) xor (A(75) and B(80)) xor (A(76) and B(79)) xor (A(77) and B(78)) xor (A(78) and B(77)) xor (A(79) and B(76)) xor (A(80) and B(75)) xor (A(81) and B(74)) xor (A(82) and B(73)) xor (A(83) and B(72)) xor (A(84) and B(71)) xor (A(85) and B(70)) xor (A(86) and B(69)) xor (A(87) and B(68)) xor (A(88) and B(67)) xor (A(89) and B(66)) xor (A(90) and B(65)) xor (A(91) and B(64)) xor (A(92) and B(63)) xor (A(93) and B(62)) xor (A(94) and B(61)) xor (A(95) and B(60)) xor (A(96) and B(59)) xor (A(97) and B(58)) xor (A(98) and B(57)) xor (A(99) and B(56)) xor (A(100) and B(55)) xor (A(101) and B(54)) xor (A(102) and B(53)) xor (A(103) and B(52)) xor (A(104) and B(51)) xor (A(105) and B(50)) xor (A(106) and B(49)) xor (A(107) and B(48)) xor (A(108) and B(47)) xor (A(109) and B(46)) xor (A(110) and B(45)) xor (A(111) and B(44)) xor (A(112) and B(43)) xor (A(113) and B(42)) xor (A(114) and B(41)) xor (A(115) and B(40)) xor (A(116) and B(39)) xor (A(117) and B(38)) xor (A(118) and B(37)) xor (A(119) and B(36)) xor (A(120) and B(35)) xor (A(121) and B(34)) xor (A(122) and B(33)) xor (A(123) and B(32)) xor (A(124) and B(31)) xor (A(125) and B(30)) xor (A(126) and B(29)) xor (A(29) and B(127)) xor (A(30) and B(126)) xor (A(31) and B(125)) xor (A(32) and B(124)) xor (A(33) and B(123)) xor (A(34) and B(122)) xor (A(35) and B(121)) xor (A(36) and B(120)) xor (A(37) and B(119)) xor (A(38) and B(118)) xor (A(39) and B(117)) xor (A(40) and B(116)) xor (A(41) and B(115)) xor (A(42) and B(114)) xor (A(43) and B(113)) xor (A(44) and B(112)) xor (A(45) and B(111)) xor (A(46) and B(110)) xor (A(47) and B(109)) xor (A(48) and B(108)) xor (A(49) and B(107)) xor (A(50) and B(106)) xor (A(51) and B(105)) xor (A(52) and B(104)) xor (A(53) and B(103)) xor (A(54) and B(102)) xor (A(55) and B(101)) xor (A(56) and B(100)) xor (A(57) and B(99)) xor (A(58) and B(98)) xor (A(59) and B(97)) xor (A(60) and B(96)) xor (A(61) and B(95)) xor (A(62) and B(94)) xor (A(63) and B(93)) xor (A(64) and B(92)) xor (A(65) and B(91)) xor (A(66) and B(90)) xor (A(67) and B(89)) xor (A(68) and B(88)) xor (A(69) and B(87)) xor (A(70) and B(86)) xor (A(71) and B(85)) xor (A(72) and B(84)) xor (A(73) and B(83)) xor (A(74) and B(82)) xor (A(75) and B(81)) xor (A(76) and B(80)) xor (A(77) and B(79)) xor (A(78) and B(78)) xor (A(79) and B(77)) xor (A(80) and B(76)) xor (A(81) and B(75)) xor (A(82) and B(74)) xor (A(83) and B(73)) xor (A(84) and B(72)) xor (A(85) and B(71)) xor (A(86) and B(70)) xor (A(87) and B(69)) xor (A(88) and B(68)) xor (A(89) and B(67)) xor (A(90) and B(66)) xor (A(91) and B(65)) xor (A(92) and B(64)) xor (A(93) and B(63)) xor (A(94) and B(62)) xor (A(95) and B(61)) xor (A(96) and B(60)) xor (A(97) and B(59)) xor (A(98) and B(58)) xor (A(99) and B(57)) xor (A(100) and B(56)) xor (A(101) and B(55)) xor (A(102) and B(54)) xor (A(103) and B(53)) xor (A(104) and B(52)) xor (A(105) and B(51)) xor (A(106) and B(50)) xor (A(107) and B(49)) xor (A(108) and B(48)) xor (A(109) and B(47)) xor (A(110) and B(46)) xor (A(111) and B(45)) xor (A(112) and B(44)) xor (A(113) and B(43)) xor (A(114) and B(42)) xor (A(115) and B(41)) xor (A(116) and B(40)) xor (A(117) and B(39)) xor (A(118) and B(38)) xor (A(119) and B(37)) xor (A(120) and B(36)) xor (A(121) and B(35)) xor (A(122) and B(34)) xor (A(123) and B(33)) xor (A(124) and B(32)) xor (A(125) and B(31)) xor (A(126) and B(30)) xor (A(30) and B(127)) xor (A(31) and B(126)) xor (A(32) and B(125)) xor (A(33) and B(124)) xor (A(34) and B(123)) xor (A(35) and B(122)) xor (A(36) and B(121)) xor (A(37) and B(120)) xor (A(38) and B(119)) xor (A(39) and B(118)) xor (A(40) and B(117)) xor (A(41) and B(116)) xor (A(42) and B(115)) xor (A(43) and B(114)) xor (A(44) and B(113)) xor (A(45) and B(112)) xor (A(46) and B(111)) xor (A(47) and B(110)) xor (A(48) and B(109)) xor (A(49) and B(108)) xor (A(50) and B(107)) xor (A(51) and B(106)) xor (A(52) and B(105)) xor (A(53) and B(104)) xor (A(54) and B(103)) xor (A(55) and B(102)) xor (A(56) and B(101)) xor (A(57) and B(100)) xor (A(58) and B(99)) xor (A(59) and B(98)) xor (A(60) and B(97)) xor (A(61) and B(96)) xor (A(62) and B(95)) xor (A(63) and B(94)) xor (A(64) and B(93)) xor (A(65) and B(92)) xor (A(66) and B(91)) xor (A(67) and B(90)) xor (A(68) and B(89)) xor (A(69) and B(88)) xor (A(70) and B(87)) xor (A(71) and B(86)) xor (A(72) and B(85)) xor (A(73) and B(84)) xor (A(74) and B(83)) xor (A(75) and B(82)) xor (A(76) and B(81)) xor (A(77) and B(80)) xor (A(78) and B(79)) xor (A(79) and B(78)) xor (A(80) and B(77)) xor (A(81) and B(76)) xor (A(82) and B(75)) xor (A(83) and B(74)) xor (A(84) and B(73)) xor (A(85) and B(72)) xor (A(86) and B(71)) xor (A(87) and B(70)) xor (A(88) and B(69)) xor (A(89) and B(68)) xor (A(90) and B(67)) xor (A(91) and B(66)) xor (A(92) and B(65)) xor (A(93) and B(64)) xor (A(94) and B(63)) xor (A(95) and B(62)) xor (A(96) and B(61)) xor (A(97) and B(60)) xor (A(98) and B(59)) xor (A(99) and B(58)) xor (A(100) and B(57)) xor (A(101) and B(56)) xor (A(102) and B(55)) xor (A(103) and B(54)) xor (A(104) and B(53)) xor (A(105) and B(52)) xor (A(106) and B(51)) xor (A(107) and B(50)) xor (A(108) and B(49)) xor (A(109) and B(48)) xor (A(110) and B(47)) xor (A(111) and B(46)) xor (A(112) and B(45)) xor (A(113) and B(44)) xor (A(114) and B(43)) xor (A(115) and B(42)) xor (A(116) and B(41)) xor (A(117) and B(40)) xor (A(118) and B(39)) xor (A(119) and B(38)) xor (A(120) and B(37)) xor (A(121) and B(36)) xor (A(122) and B(35)) xor (A(123) and B(34)) xor (A(124) and B(33)) xor (A(125) and B(32)) xor (A(126) and B(32));
    C(31)  <= (A(0) and B(31)) xor (A(1) and B(30)) xor (A(2) and B(29)) xor (A(3) and B(28)) xor (A(4) and B(27)) xor (A(5) and B(26)) xor (A(6) and B(25)) xor (A(7) and B(24)) xor (A(8) and B(23)) xor (A(9) and B(23)) xor (A(10) and B(21)) xor (A(11) and B(20)) xor (A(12) and B(19)) xor (A(13) and B(18)) xor (A(14) and B(17)) xor (A(15) and B(16)) xor (A(16) and B(15)) xor (A(17) and B(14)) xor (A(18) and B(13)) xor (A(19) and B(12)) xor (A(20) and B(11)) xor (A(21) and B(10)) xor (A(23) and B(9)) xor (A(23) and B(8)) xor (A(24) and B(7)) xor (A(25) and B(6)) xor (A(26) and B(5)) xor (A(27) and B(4)) xor (A(28) and B(3)) xor (A(29) and B(2)) xor (A(30) and B(1)) xor (A(31) and B(0)) xor (A(24) and B(127)) xor (A(25) and B(126)) xor (A(26) and B(125)) xor (A(27) and B(124)) xor (A(28) and B(123)) xor (A(29) and B(122)) xor (A(30) and B(121)) xor (A(31) and B(120)) xor (A(32) and B(119)) xor (A(33) and B(118)) xor (A(34) and B(117)) xor (A(35) and B(116)) xor (A(36) and B(115)) xor (A(37) and B(114)) xor (A(38) and B(113)) xor (A(39) and B(112)) xor (A(40) and B(111)) xor (A(41) and B(110)) xor (A(42) and B(109)) xor (A(43) and B(108)) xor (A(44) and B(107)) xor (A(45) and B(106)) xor (A(46) and B(105)) xor (A(47) and B(104)) xor (A(48) and B(103)) xor (A(49) and B(102)) xor (A(50) and B(101)) xor (A(51) and B(100)) xor (A(52) and B(99)) xor (A(53) and B(98)) xor (A(54) and B(97)) xor (A(55) and B(96)) xor (A(56) and B(95)) xor (A(57) and B(94)) xor (A(58) and B(93)) xor (A(59) and B(92)) xor (A(60) and B(91)) xor (A(61) and B(90)) xor (A(62) and B(89)) xor (A(63) and B(88)) xor (A(64) and B(87)) xor (A(65) and B(86)) xor (A(66) and B(85)) xor (A(67) and B(84)) xor (A(68) and B(83)) xor (A(69) and B(82)) xor (A(70) and B(81)) xor (A(71) and B(80)) xor (A(72) and B(79)) xor (A(73) and B(78)) xor (A(74) and B(77)) xor (A(75) and B(76)) xor (A(76) and B(75)) xor (A(77) and B(74)) xor (A(78) and B(73)) xor (A(79) and B(72)) xor (A(80) and B(71)) xor (A(81) and B(70)) xor (A(82) and B(69)) xor (A(83) and B(68)) xor (A(84) and B(67)) xor (A(85) and B(66)) xor (A(86) and B(65)) xor (A(87) and B(64)) xor (A(88) and B(63)) xor (A(89) and B(62)) xor (A(90) and B(61)) xor (A(91) and B(60)) xor (A(92) and B(59)) xor (A(93) and B(58)) xor (A(94) and B(57)) xor (A(95) and B(56)) xor (A(96) and B(55)) xor (A(97) and B(54)) xor (A(98) and B(53)) xor (A(99) and B(52)) xor (A(100) and B(51)) xor (A(101) and B(50)) xor (A(102) and B(49)) xor (A(103) and B(48)) xor (A(104) and B(47)) xor (A(105) and B(46)) xor (A(106) and B(45)) xor (A(107) and B(44)) xor (A(108) and B(43)) xor (A(109) and B(42)) xor (A(110) and B(41)) xor (A(111) and B(40)) xor (A(112) and B(39)) xor (A(113) and B(38)) xor (A(114) and B(37)) xor (A(115) and B(36)) xor (A(116) and B(35)) xor (A(117) and B(34)) xor (A(118) and B(33)) xor (A(119) and B(32)) xor (A(120) and B(31)) xor (A(121) and B(30)) xor (A(122) and B(29)) xor (A(123) and B(28)) xor (A(124) and B(27)) xor (A(125) and B(26)) xor (A(126) and B(25)) xor (A(29) and B(127)) xor (A(30) and B(126)) xor (A(31) and B(125)) xor (A(32) and B(124)) xor (A(33) and B(123)) xor (A(34) and B(122)) xor (A(35) and B(121)) xor (A(36) and B(120)) xor (A(37) and B(119)) xor (A(38) and B(118)) xor (A(39) and B(117)) xor (A(40) and B(116)) xor (A(41) and B(115)) xor (A(42) and B(114)) xor (A(43) and B(113)) xor (A(44) and B(112)) xor (A(45) and B(111)) xor (A(46) and B(110)) xor (A(47) and B(109)) xor (A(48) and B(108)) xor (A(49) and B(107)) xor (A(50) and B(106)) xor (A(51) and B(105)) xor (A(52) and B(104)) xor (A(53) and B(103)) xor (A(54) and B(102)) xor (A(55) and B(101)) xor (A(56) and B(100)) xor (A(57) and B(99)) xor (A(58) and B(98)) xor (A(59) and B(97)) xor (A(60) and B(96)) xor (A(61) and B(95)) xor (A(62) and B(94)) xor (A(63) and B(93)) xor (A(64) and B(92)) xor (A(65) and B(91)) xor (A(66) and B(90)) xor (A(67) and B(89)) xor (A(68) and B(88)) xor (A(69) and B(87)) xor (A(70) and B(86)) xor (A(71) and B(85)) xor (A(72) and B(84)) xor (A(73) and B(83)) xor (A(74) and B(82)) xor (A(75) and B(81)) xor (A(76) and B(80)) xor (A(77) and B(79)) xor (A(78) and B(78)) xor (A(79) and B(77)) xor (A(80) and B(76)) xor (A(81) and B(75)) xor (A(82) and B(74)) xor (A(83) and B(73)) xor (A(84) and B(72)) xor (A(85) and B(71)) xor (A(86) and B(70)) xor (A(87) and B(69)) xor (A(88) and B(68)) xor (A(89) and B(67)) xor (A(90) and B(66)) xor (A(91) and B(65)) xor (A(92) and B(64)) xor (A(93) and B(63)) xor (A(94) and B(62)) xor (A(95) and B(61)) xor (A(96) and B(60)) xor (A(97) and B(59)) xor (A(98) and B(58)) xor (A(99) and B(57)) xor (A(100) and B(56)) xor (A(101) and B(55)) xor (A(102) and B(54)) xor (A(103) and B(53)) xor (A(104) and B(52)) xor (A(105) and B(51)) xor (A(106) and B(50)) xor (A(107) and B(49)) xor (A(108) and B(48)) xor (A(109) and B(47)) xor (A(110) and B(46)) xor (A(111) and B(45)) xor (A(112) and B(44)) xor (A(113) and B(43)) xor (A(114) and B(42)) xor (A(115) and B(41)) xor (A(116) and B(40)) xor (A(117) and B(39)) xor (A(118) and B(38)) xor (A(119) and B(37)) xor (A(120) and B(36)) xor (A(121) and B(35)) xor (A(122) and B(34)) xor (A(123) and B(33)) xor (A(124) and B(32)) xor (A(125) and B(31)) xor (A(126) and B(30)) xor (A(30) and B(127)) xor (A(31) and B(126)) xor (A(32) and B(125)) xor (A(33) and B(124)) xor (A(34) and B(123)) xor (A(35) and B(122)) xor (A(36) and B(121)) xor (A(37) and B(120)) xor (A(38) and B(119)) xor (A(39) and B(118)) xor (A(40) and B(117)) xor (A(41) and B(116)) xor (A(42) and B(115)) xor (A(43) and B(114)) xor (A(44) and B(113)) xor (A(45) and B(112)) xor (A(46) and B(111)) xor (A(47) and B(110)) xor (A(48) and B(109)) xor (A(49) and B(108)) xor (A(50) and B(107)) xor (A(51) and B(106)) xor (A(52) and B(105)) xor (A(53) and B(104)) xor (A(54) and B(103)) xor (A(55) and B(102)) xor (A(56) and B(101)) xor (A(57) and B(100)) xor (A(58) and B(99)) xor (A(59) and B(98)) xor (A(60) and B(97)) xor (A(61) and B(96)) xor (A(62) and B(95)) xor (A(63) and B(94)) xor (A(64) and B(93)) xor (A(65) and B(92)) xor (A(66) and B(91)) xor (A(67) and B(90)) xor (A(68) and B(89)) xor (A(69) and B(88)) xor (A(70) and B(87)) xor (A(71) and B(86)) xor (A(72) and B(85)) xor (A(73) and B(84)) xor (A(74) and B(83)) xor (A(75) and B(82)) xor (A(76) and B(81)) xor (A(77) and B(80)) xor (A(78) and B(79)) xor (A(79) and B(78)) xor (A(80) and B(77)) xor (A(81) and B(76)) xor (A(82) and B(75)) xor (A(83) and B(74)) xor (A(84) and B(73)) xor (A(85) and B(72)) xor (A(86) and B(71)) xor (A(87) and B(70)) xor (A(88) and B(69)) xor (A(89) and B(68)) xor (A(90) and B(67)) xor (A(91) and B(66)) xor (A(92) and B(65)) xor (A(93) and B(64)) xor (A(94) and B(63)) xor (A(95) and B(62)) xor (A(96) and B(61)) xor (A(97) and B(60)) xor (A(98) and B(59)) xor (A(99) and B(58)) xor (A(100) and B(57)) xor (A(101) and B(56)) xor (A(102) and B(55)) xor (A(103) and B(54)) xor (A(104) and B(53)) xor (A(105) and B(52)) xor (A(106) and B(51)) xor (A(107) and B(50)) xor (A(108) and B(49)) xor (A(109) and B(48)) xor (A(110) and B(47)) xor (A(111) and B(46)) xor (A(112) and B(45)) xor (A(113) and B(44)) xor (A(114) and B(43)) xor (A(115) and B(42)) xor (A(116) and B(41)) xor (A(117) and B(40)) xor (A(118) and B(39)) xor (A(119) and B(38)) xor (A(120) and B(37)) xor (A(121) and B(36)) xor (A(122) and B(35)) xor (A(123) and B(34)) xor (A(124) and B(33)) xor (A(125) and B(32)) xor (A(126) and B(31)) xor (A(31) and B(127)) xor (A(32) and B(126)) xor (A(33) and B(125)) xor (A(34) and B(124)) xor (A(35) and B(123)) xor (A(36) and B(122)) xor (A(37) and B(121)) xor (A(38) and B(120)) xor (A(39) and B(119)) xor (A(40) and B(118)) xor (A(41) and B(117)) xor (A(42) and B(116)) xor (A(43) and B(115)) xor (A(44) and B(114)) xor (A(45) and B(113)) xor (A(46) and B(112)) xor (A(47) and B(111)) xor (A(48) and B(110)) xor (A(49) and B(109)) xor (A(50) and B(108)) xor (A(51) and B(107)) xor (A(52) and B(106)) xor (A(53) and B(105)) xor (A(54) and B(104)) xor (A(55) and B(103)) xor (A(56) and B(102)) xor (A(57) and B(101)) xor (A(58) and B(100)) xor (A(59) and B(99)) xor (A(60) and B(98)) xor (A(61) and B(97)) xor (A(62) and B(96)) xor (A(63) and B(95)) xor (A(64) and B(94)) xor (A(65) and B(93)) xor (A(66) and B(92)) xor (A(67) and B(91)) xor (A(68) and B(90)) xor (A(69) and B(89)) xor (A(70) and B(88)) xor (A(71) and B(87)) xor (A(72) and B(86)) xor (A(73) and B(85)) xor (A(74) and B(84)) xor (A(75) and B(83)) xor (A(76) and B(82)) xor (A(77) and B(81)) xor (A(78) and B(80)) xor (A(79) and B(79)) xor (A(80) and B(78)) xor (A(81) and B(77)) xor (A(82) and B(76)) xor (A(83) and B(75)) xor (A(84) and B(74)) xor (A(85) and B(73)) xor (A(86) and B(72)) xor (A(87) and B(71)) xor (A(88) and B(70)) xor (A(89) and B(69)) xor (A(90) and B(68)) xor (A(91) and B(67)) xor (A(92) and B(66)) xor (A(93) and B(65)) xor (A(94) and B(64)) xor (A(95) and B(63)) xor (A(96) and B(62)) xor (A(97) and B(61)) xor (A(98) and B(60)) xor (A(99) and B(59)) xor (A(100) and B(58)) xor (A(101) and B(57)) xor (A(102) and B(56)) xor (A(103) and B(55)) xor (A(104) and B(54)) xor (A(105) and B(53)) xor (A(106) and B(52)) xor (A(107) and B(51)) xor (A(108) and B(50)) xor (A(109) and B(49)) xor (A(110) and B(48)) xor (A(111) and B(47)) xor (A(112) and B(46)) xor (A(113) and B(45)) xor (A(114) and B(44)) xor (A(115) and B(43)) xor (A(116) and B(42)) xor (A(117) and B(41)) xor (A(118) and B(40)) xor (A(119) and B(39)) xor (A(120) and B(38)) xor (A(121) and B(37)) xor (A(122) and B(36)) xor (A(123) and B(35)) xor (A(124) and B(34)) xor (A(125) and B(33)) xor (A(126) and B(33));
    C(32)  <= (A(0) and B(32)) xor (A(1) and B(31)) xor (A(2) and B(30)) xor (A(3) and B(29)) xor (A(4) and B(28)) xor (A(5) and B(27)) xor (A(6) and B(26)) xor (A(7) and B(25)) xor (A(8) and B(24)) xor (A(9) and B(23)) xor (A(10) and B(23)) xor (A(11) and B(21)) xor (A(12) and B(20)) xor (A(13) and B(19)) xor (A(14) and B(18)) xor (A(15) and B(17)) xor (A(16) and B(16)) xor (A(17) and B(15)) xor (A(18) and B(14)) xor (A(19) and B(13)) xor (A(20) and B(12)) xor (A(21) and B(11)) xor (A(23) and B(10)) xor (A(23) and B(9)) xor (A(24) and B(8)) xor (A(25) and B(7)) xor (A(26) and B(6)) xor (A(27) and B(5)) xor (A(28) and B(4)) xor (A(29) and B(3)) xor (A(30) and B(2)) xor (A(31) and B(1)) xor (A(32) and B(0)) xor (A(25) and B(127)) xor (A(26) and B(126)) xor (A(27) and B(125)) xor (A(28) and B(124)) xor (A(29) and B(123)) xor (A(30) and B(122)) xor (A(31) and B(121)) xor (A(32) and B(120)) xor (A(33) and B(119)) xor (A(34) and B(118)) xor (A(35) and B(117)) xor (A(36) and B(116)) xor (A(37) and B(115)) xor (A(38) and B(114)) xor (A(39) and B(113)) xor (A(40) and B(112)) xor (A(41) and B(111)) xor (A(42) and B(110)) xor (A(43) and B(109)) xor (A(44) and B(108)) xor (A(45) and B(107)) xor (A(46) and B(106)) xor (A(47) and B(105)) xor (A(48) and B(104)) xor (A(49) and B(103)) xor (A(50) and B(102)) xor (A(51) and B(101)) xor (A(52) and B(100)) xor (A(53) and B(99)) xor (A(54) and B(98)) xor (A(55) and B(97)) xor (A(56) and B(96)) xor (A(57) and B(95)) xor (A(58) and B(94)) xor (A(59) and B(93)) xor (A(60) and B(92)) xor (A(61) and B(91)) xor (A(62) and B(90)) xor (A(63) and B(89)) xor (A(64) and B(88)) xor (A(65) and B(87)) xor (A(66) and B(86)) xor (A(67) and B(85)) xor (A(68) and B(84)) xor (A(69) and B(83)) xor (A(70) and B(82)) xor (A(71) and B(81)) xor (A(72) and B(80)) xor (A(73) and B(79)) xor (A(74) and B(78)) xor (A(75) and B(77)) xor (A(76) and B(76)) xor (A(77) and B(75)) xor (A(78) and B(74)) xor (A(79) and B(73)) xor (A(80) and B(72)) xor (A(81) and B(71)) xor (A(82) and B(70)) xor (A(83) and B(69)) xor (A(84) and B(68)) xor (A(85) and B(67)) xor (A(86) and B(66)) xor (A(87) and B(65)) xor (A(88) and B(64)) xor (A(89) and B(63)) xor (A(90) and B(62)) xor (A(91) and B(61)) xor (A(92) and B(60)) xor (A(93) and B(59)) xor (A(94) and B(58)) xor (A(95) and B(57)) xor (A(96) and B(56)) xor (A(97) and B(55)) xor (A(98) and B(54)) xor (A(99) and B(53)) xor (A(100) and B(52)) xor (A(101) and B(51)) xor (A(102) and B(50)) xor (A(103) and B(49)) xor (A(104) and B(48)) xor (A(105) and B(47)) xor (A(106) and B(46)) xor (A(107) and B(45)) xor (A(108) and B(44)) xor (A(109) and B(43)) xor (A(110) and B(42)) xor (A(111) and B(41)) xor (A(112) and B(40)) xor (A(113) and B(39)) xor (A(114) and B(38)) xor (A(115) and B(37)) xor (A(116) and B(36)) xor (A(117) and B(35)) xor (A(118) and B(34)) xor (A(119) and B(33)) xor (A(120) and B(32)) xor (A(121) and B(31)) xor (A(122) and B(30)) xor (A(123) and B(29)) xor (A(124) and B(28)) xor (A(125) and B(27)) xor (A(126) and B(26)) xor (A(30) and B(127)) xor (A(31) and B(126)) xor (A(32) and B(125)) xor (A(33) and B(124)) xor (A(34) and B(123)) xor (A(35) and B(122)) xor (A(36) and B(121)) xor (A(37) and B(120)) xor (A(38) and B(119)) xor (A(39) and B(118)) xor (A(40) and B(117)) xor (A(41) and B(116)) xor (A(42) and B(115)) xor (A(43) and B(114)) xor (A(44) and B(113)) xor (A(45) and B(112)) xor (A(46) and B(111)) xor (A(47) and B(110)) xor (A(48) and B(109)) xor (A(49) and B(108)) xor (A(50) and B(107)) xor (A(51) and B(106)) xor (A(52) and B(105)) xor (A(53) and B(104)) xor (A(54) and B(103)) xor (A(55) and B(102)) xor (A(56) and B(101)) xor (A(57) and B(100)) xor (A(58) and B(99)) xor (A(59) and B(98)) xor (A(60) and B(97)) xor (A(61) and B(96)) xor (A(62) and B(95)) xor (A(63) and B(94)) xor (A(64) and B(93)) xor (A(65) and B(92)) xor (A(66) and B(91)) xor (A(67) and B(90)) xor (A(68) and B(89)) xor (A(69) and B(88)) xor (A(70) and B(87)) xor (A(71) and B(86)) xor (A(72) and B(85)) xor (A(73) and B(84)) xor (A(74) and B(83)) xor (A(75) and B(82)) xor (A(76) and B(81)) xor (A(77) and B(80)) xor (A(78) and B(79)) xor (A(79) and B(78)) xor (A(80) and B(77)) xor (A(81) and B(76)) xor (A(82) and B(75)) xor (A(83) and B(74)) xor (A(84) and B(73)) xor (A(85) and B(72)) xor (A(86) and B(71)) xor (A(87) and B(70)) xor (A(88) and B(69)) xor (A(89) and B(68)) xor (A(90) and B(67)) xor (A(91) and B(66)) xor (A(92) and B(65)) xor (A(93) and B(64)) xor (A(94) and B(63)) xor (A(95) and B(62)) xor (A(96) and B(61)) xor (A(97) and B(60)) xor (A(98) and B(59)) xor (A(99) and B(58)) xor (A(100) and B(57)) xor (A(101) and B(56)) xor (A(102) and B(55)) xor (A(103) and B(54)) xor (A(104) and B(53)) xor (A(105) and B(52)) xor (A(106) and B(51)) xor (A(107) and B(50)) xor (A(108) and B(49)) xor (A(109) and B(48)) xor (A(110) and B(47)) xor (A(111) and B(46)) xor (A(112) and B(45)) xor (A(113) and B(44)) xor (A(114) and B(43)) xor (A(115) and B(42)) xor (A(116) and B(41)) xor (A(117) and B(40)) xor (A(118) and B(39)) xor (A(119) and B(38)) xor (A(120) and B(37)) xor (A(121) and B(36)) xor (A(122) and B(35)) xor (A(123) and B(34)) xor (A(124) and B(33)) xor (A(125) and B(32)) xor (A(126) and B(31)) xor (A(31) and B(127)) xor (A(32) and B(126)) xor (A(33) and B(125)) xor (A(34) and B(124)) xor (A(35) and B(123)) xor (A(36) and B(122)) xor (A(37) and B(121)) xor (A(38) and B(120)) xor (A(39) and B(119)) xor (A(40) and B(118)) xor (A(41) and B(117)) xor (A(42) and B(116)) xor (A(43) and B(115)) xor (A(44) and B(114)) xor (A(45) and B(113)) xor (A(46) and B(112)) xor (A(47) and B(111)) xor (A(48) and B(110)) xor (A(49) and B(109)) xor (A(50) and B(108)) xor (A(51) and B(107)) xor (A(52) and B(106)) xor (A(53) and B(105)) xor (A(54) and B(104)) xor (A(55) and B(103)) xor (A(56) and B(102)) xor (A(57) and B(101)) xor (A(58) and B(100)) xor (A(59) and B(99)) xor (A(60) and B(98)) xor (A(61) and B(97)) xor (A(62) and B(96)) xor (A(63) and B(95)) xor (A(64) and B(94)) xor (A(65) and B(93)) xor (A(66) and B(92)) xor (A(67) and B(91)) xor (A(68) and B(90)) xor (A(69) and B(89)) xor (A(70) and B(88)) xor (A(71) and B(87)) xor (A(72) and B(86)) xor (A(73) and B(85)) xor (A(74) and B(84)) xor (A(75) and B(83)) xor (A(76) and B(82)) xor (A(77) and B(81)) xor (A(78) and B(80)) xor (A(79) and B(79)) xor (A(80) and B(78)) xor (A(81) and B(77)) xor (A(82) and B(76)) xor (A(83) and B(75)) xor (A(84) and B(74)) xor (A(85) and B(73)) xor (A(86) and B(72)) xor (A(87) and B(71)) xor (A(88) and B(70)) xor (A(89) and B(69)) xor (A(90) and B(68)) xor (A(91) and B(67)) xor (A(92) and B(66)) xor (A(93) and B(65)) xor (A(94) and B(64)) xor (A(95) and B(63)) xor (A(96) and B(62)) xor (A(97) and B(61)) xor (A(98) and B(60)) xor (A(99) and B(59)) xor (A(100) and B(58)) xor (A(101) and B(57)) xor (A(102) and B(56)) xor (A(103) and B(55)) xor (A(104) and B(54)) xor (A(105) and B(53)) xor (A(106) and B(52)) xor (A(107) and B(51)) xor (A(108) and B(50)) xor (A(109) and B(49)) xor (A(110) and B(48)) xor (A(111) and B(47)) xor (A(112) and B(46)) xor (A(113) and B(45)) xor (A(114) and B(44)) xor (A(115) and B(43)) xor (A(116) and B(42)) xor (A(117) and B(41)) xor (A(118) and B(40)) xor (A(119) and B(39)) xor (A(120) and B(38)) xor (A(121) and B(37)) xor (A(122) and B(36)) xor (A(123) and B(35)) xor (A(124) and B(34)) xor (A(125) and B(33)) xor (A(126) and B(32)) xor (A(32) and B(127)) xor (A(33) and B(126)) xor (A(34) and B(125)) xor (A(35) and B(124)) xor (A(36) and B(123)) xor (A(37) and B(122)) xor (A(38) and B(121)) xor (A(39) and B(120)) xor (A(40) and B(119)) xor (A(41) and B(118)) xor (A(42) and B(117)) xor (A(43) and B(116)) xor (A(44) and B(115)) xor (A(45) and B(114)) xor (A(46) and B(113)) xor (A(47) and B(112)) xor (A(48) and B(111)) xor (A(49) and B(110)) xor (A(50) and B(109)) xor (A(51) and B(108)) xor (A(52) and B(107)) xor (A(53) and B(106)) xor (A(54) and B(105)) xor (A(55) and B(104)) xor (A(56) and B(103)) xor (A(57) and B(102)) xor (A(58) and B(101)) xor (A(59) and B(100)) xor (A(60) and B(99)) xor (A(61) and B(98)) xor (A(62) and B(97)) xor (A(63) and B(96)) xor (A(64) and B(95)) xor (A(65) and B(94)) xor (A(66) and B(93)) xor (A(67) and B(92)) xor (A(68) and B(91)) xor (A(69) and B(90)) xor (A(70) and B(89)) xor (A(71) and B(88)) xor (A(72) and B(87)) xor (A(73) and B(86)) xor (A(74) and B(85)) xor (A(75) and B(84)) xor (A(76) and B(83)) xor (A(77) and B(82)) xor (A(78) and B(81)) xor (A(79) and B(80)) xor (A(80) and B(79)) xor (A(81) and B(78)) xor (A(82) and B(77)) xor (A(83) and B(76)) xor (A(84) and B(75)) xor (A(85) and B(74)) xor (A(86) and B(73)) xor (A(87) and B(72)) xor (A(88) and B(71)) xor (A(89) and B(70)) xor (A(90) and B(69)) xor (A(91) and B(68)) xor (A(92) and B(67)) xor (A(93) and B(66)) xor (A(94) and B(65)) xor (A(95) and B(64)) xor (A(96) and B(63)) xor (A(97) and B(62)) xor (A(98) and B(61)) xor (A(99) and B(60)) xor (A(100) and B(59)) xor (A(101) and B(58)) xor (A(102) and B(57)) xor (A(103) and B(56)) xor (A(104) and B(55)) xor (A(105) and B(54)) xor (A(106) and B(53)) xor (A(107) and B(52)) xor (A(108) and B(51)) xor (A(109) and B(50)) xor (A(110) and B(49)) xor (A(111) and B(48)) xor (A(112) and B(47)) xor (A(113) and B(46)) xor (A(114) and B(45)) xor (A(115) and B(44)) xor (A(116) and B(43)) xor (A(117) and B(42)) xor (A(118) and B(41)) xor (A(119) and B(40)) xor (A(120) and B(39)) xor (A(121) and B(38)) xor (A(122) and B(37)) xor (A(123) and B(36)) xor (A(124) and B(35)) xor (A(125) and B(34)) xor (A(126) and B(34));
    C(33)  <= (A(0) and B(33)) xor (A(1) and B(32)) xor (A(2) and B(31)) xor (A(3) and B(30)) xor (A(4) and B(29)) xor (A(5) and B(28)) xor (A(6) and B(27)) xor (A(7) and B(26)) xor (A(8) and B(25)) xor (A(9) and B(24)) xor (A(10) and B(23)) xor (A(11) and B(23)) xor (A(12) and B(21)) xor (A(13) and B(20)) xor (A(14) and B(19)) xor (A(15) and B(18)) xor (A(16) and B(17)) xor (A(17) and B(16)) xor (A(18) and B(15)) xor (A(19) and B(14)) xor (A(20) and B(13)) xor (A(21) and B(12)) xor (A(23) and B(11)) xor (A(23) and B(10)) xor (A(24) and B(9)) xor (A(25) and B(8)) xor (A(26) and B(7)) xor (A(27) and B(6)) xor (A(28) and B(5)) xor (A(29) and B(4)) xor (A(30) and B(3)) xor (A(31) and B(2)) xor (A(32) and B(1)) xor (A(33) and B(0)) xor (A(26) and B(127)) xor (A(27) and B(126)) xor (A(28) and B(125)) xor (A(29) and B(124)) xor (A(30) and B(123)) xor (A(31) and B(122)) xor (A(32) and B(121)) xor (A(33) and B(120)) xor (A(34) and B(119)) xor (A(35) and B(118)) xor (A(36) and B(117)) xor (A(37) and B(116)) xor (A(38) and B(115)) xor (A(39) and B(114)) xor (A(40) and B(113)) xor (A(41) and B(112)) xor (A(42) and B(111)) xor (A(43) and B(110)) xor (A(44) and B(109)) xor (A(45) and B(108)) xor (A(46) and B(107)) xor (A(47) and B(106)) xor (A(48) and B(105)) xor (A(49) and B(104)) xor (A(50) and B(103)) xor (A(51) and B(102)) xor (A(52) and B(101)) xor (A(53) and B(100)) xor (A(54) and B(99)) xor (A(55) and B(98)) xor (A(56) and B(97)) xor (A(57) and B(96)) xor (A(58) and B(95)) xor (A(59) and B(94)) xor (A(60) and B(93)) xor (A(61) and B(92)) xor (A(62) and B(91)) xor (A(63) and B(90)) xor (A(64) and B(89)) xor (A(65) and B(88)) xor (A(66) and B(87)) xor (A(67) and B(86)) xor (A(68) and B(85)) xor (A(69) and B(84)) xor (A(70) and B(83)) xor (A(71) and B(82)) xor (A(72) and B(81)) xor (A(73) and B(80)) xor (A(74) and B(79)) xor (A(75) and B(78)) xor (A(76) and B(77)) xor (A(77) and B(76)) xor (A(78) and B(75)) xor (A(79) and B(74)) xor (A(80) and B(73)) xor (A(81) and B(72)) xor (A(82) and B(71)) xor (A(83) and B(70)) xor (A(84) and B(69)) xor (A(85) and B(68)) xor (A(86) and B(67)) xor (A(87) and B(66)) xor (A(88) and B(65)) xor (A(89) and B(64)) xor (A(90) and B(63)) xor (A(91) and B(62)) xor (A(92) and B(61)) xor (A(93) and B(60)) xor (A(94) and B(59)) xor (A(95) and B(58)) xor (A(96) and B(57)) xor (A(97) and B(56)) xor (A(98) and B(55)) xor (A(99) and B(54)) xor (A(100) and B(53)) xor (A(101) and B(52)) xor (A(102) and B(51)) xor (A(103) and B(50)) xor (A(104) and B(49)) xor (A(105) and B(48)) xor (A(106) and B(47)) xor (A(107) and B(46)) xor (A(108) and B(45)) xor (A(109) and B(44)) xor (A(110) and B(43)) xor (A(111) and B(42)) xor (A(112) and B(41)) xor (A(113) and B(40)) xor (A(114) and B(39)) xor (A(115) and B(38)) xor (A(116) and B(37)) xor (A(117) and B(36)) xor (A(118) and B(35)) xor (A(119) and B(34)) xor (A(120) and B(33)) xor (A(121) and B(32)) xor (A(122) and B(31)) xor (A(123) and B(30)) xor (A(124) and B(29)) xor (A(125) and B(28)) xor (A(126) and B(27)) xor (A(31) and B(127)) xor (A(32) and B(126)) xor (A(33) and B(125)) xor (A(34) and B(124)) xor (A(35) and B(123)) xor (A(36) and B(122)) xor (A(37) and B(121)) xor (A(38) and B(120)) xor (A(39) and B(119)) xor (A(40) and B(118)) xor (A(41) and B(117)) xor (A(42) and B(116)) xor (A(43) and B(115)) xor (A(44) and B(114)) xor (A(45) and B(113)) xor (A(46) and B(112)) xor (A(47) and B(111)) xor (A(48) and B(110)) xor (A(49) and B(109)) xor (A(50) and B(108)) xor (A(51) and B(107)) xor (A(52) and B(106)) xor (A(53) and B(105)) xor (A(54) and B(104)) xor (A(55) and B(103)) xor (A(56) and B(102)) xor (A(57) and B(101)) xor (A(58) and B(100)) xor (A(59) and B(99)) xor (A(60) and B(98)) xor (A(61) and B(97)) xor (A(62) and B(96)) xor (A(63) and B(95)) xor (A(64) and B(94)) xor (A(65) and B(93)) xor (A(66) and B(92)) xor (A(67) and B(91)) xor (A(68) and B(90)) xor (A(69) and B(89)) xor (A(70) and B(88)) xor (A(71) and B(87)) xor (A(72) and B(86)) xor (A(73) and B(85)) xor (A(74) and B(84)) xor (A(75) and B(83)) xor (A(76) and B(82)) xor (A(77) and B(81)) xor (A(78) and B(80)) xor (A(79) and B(79)) xor (A(80) and B(78)) xor (A(81) and B(77)) xor (A(82) and B(76)) xor (A(83) and B(75)) xor (A(84) and B(74)) xor (A(85) and B(73)) xor (A(86) and B(72)) xor (A(87) and B(71)) xor (A(88) and B(70)) xor (A(89) and B(69)) xor (A(90) and B(68)) xor (A(91) and B(67)) xor (A(92) and B(66)) xor (A(93) and B(65)) xor (A(94) and B(64)) xor (A(95) and B(63)) xor (A(96) and B(62)) xor (A(97) and B(61)) xor (A(98) and B(60)) xor (A(99) and B(59)) xor (A(100) and B(58)) xor (A(101) and B(57)) xor (A(102) and B(56)) xor (A(103) and B(55)) xor (A(104) and B(54)) xor (A(105) and B(53)) xor (A(106) and B(52)) xor (A(107) and B(51)) xor (A(108) and B(50)) xor (A(109) and B(49)) xor (A(110) and B(48)) xor (A(111) and B(47)) xor (A(112) and B(46)) xor (A(113) and B(45)) xor (A(114) and B(44)) xor (A(115) and B(43)) xor (A(116) and B(42)) xor (A(117) and B(41)) xor (A(118) and B(40)) xor (A(119) and B(39)) xor (A(120) and B(38)) xor (A(121) and B(37)) xor (A(122) and B(36)) xor (A(123) and B(35)) xor (A(124) and B(34)) xor (A(125) and B(33)) xor (A(126) and B(32)) xor (A(32) and B(127)) xor (A(33) and B(126)) xor (A(34) and B(125)) xor (A(35) and B(124)) xor (A(36) and B(123)) xor (A(37) and B(122)) xor (A(38) and B(121)) xor (A(39) and B(120)) xor (A(40) and B(119)) xor (A(41) and B(118)) xor (A(42) and B(117)) xor (A(43) and B(116)) xor (A(44) and B(115)) xor (A(45) and B(114)) xor (A(46) and B(113)) xor (A(47) and B(112)) xor (A(48) and B(111)) xor (A(49) and B(110)) xor (A(50) and B(109)) xor (A(51) and B(108)) xor (A(52) and B(107)) xor (A(53) and B(106)) xor (A(54) and B(105)) xor (A(55) and B(104)) xor (A(56) and B(103)) xor (A(57) and B(102)) xor (A(58) and B(101)) xor (A(59) and B(100)) xor (A(60) and B(99)) xor (A(61) and B(98)) xor (A(62) and B(97)) xor (A(63) and B(96)) xor (A(64) and B(95)) xor (A(65) and B(94)) xor (A(66) and B(93)) xor (A(67) and B(92)) xor (A(68) and B(91)) xor (A(69) and B(90)) xor (A(70) and B(89)) xor (A(71) and B(88)) xor (A(72) and B(87)) xor (A(73) and B(86)) xor (A(74) and B(85)) xor (A(75) and B(84)) xor (A(76) and B(83)) xor (A(77) and B(82)) xor (A(78) and B(81)) xor (A(79) and B(80)) xor (A(80) and B(79)) xor (A(81) and B(78)) xor (A(82) and B(77)) xor (A(83) and B(76)) xor (A(84) and B(75)) xor (A(85) and B(74)) xor (A(86) and B(73)) xor (A(87) and B(72)) xor (A(88) and B(71)) xor (A(89) and B(70)) xor (A(90) and B(69)) xor (A(91) and B(68)) xor (A(92) and B(67)) xor (A(93) and B(66)) xor (A(94) and B(65)) xor (A(95) and B(64)) xor (A(96) and B(63)) xor (A(97) and B(62)) xor (A(98) and B(61)) xor (A(99) and B(60)) xor (A(100) and B(59)) xor (A(101) and B(58)) xor (A(102) and B(57)) xor (A(103) and B(56)) xor (A(104) and B(55)) xor (A(105) and B(54)) xor (A(106) and B(53)) xor (A(107) and B(52)) xor (A(108) and B(51)) xor (A(109) and B(50)) xor (A(110) and B(49)) xor (A(111) and B(48)) xor (A(112) and B(47)) xor (A(113) and B(46)) xor (A(114) and B(45)) xor (A(115) and B(44)) xor (A(116) and B(43)) xor (A(117) and B(42)) xor (A(118) and B(41)) xor (A(119) and B(40)) xor (A(120) and B(39)) xor (A(121) and B(38)) xor (A(122) and B(37)) xor (A(123) and B(36)) xor (A(124) and B(35)) xor (A(125) and B(34)) xor (A(126) and B(33)) xor (A(33) and B(127)) xor (A(34) and B(126)) xor (A(35) and B(125)) xor (A(36) and B(124)) xor (A(37) and B(123)) xor (A(38) and B(122)) xor (A(39) and B(121)) xor (A(40) and B(120)) xor (A(41) and B(119)) xor (A(42) and B(118)) xor (A(43) and B(117)) xor (A(44) and B(116)) xor (A(45) and B(115)) xor (A(46) and B(114)) xor (A(47) and B(113)) xor (A(48) and B(112)) xor (A(49) and B(111)) xor (A(50) and B(110)) xor (A(51) and B(109)) xor (A(52) and B(108)) xor (A(53) and B(107)) xor (A(54) and B(106)) xor (A(55) and B(105)) xor (A(56) and B(104)) xor (A(57) and B(103)) xor (A(58) and B(102)) xor (A(59) and B(101)) xor (A(60) and B(100)) xor (A(61) and B(99)) xor (A(62) and B(98)) xor (A(63) and B(97)) xor (A(64) and B(96)) xor (A(65) and B(95)) xor (A(66) and B(94)) xor (A(67) and B(93)) xor (A(68) and B(92)) xor (A(69) and B(91)) xor (A(70) and B(90)) xor (A(71) and B(89)) xor (A(72) and B(88)) xor (A(73) and B(87)) xor (A(74) and B(86)) xor (A(75) and B(85)) xor (A(76) and B(84)) xor (A(77) and B(83)) xor (A(78) and B(82)) xor (A(79) and B(81)) xor (A(80) and B(80)) xor (A(81) and B(79)) xor (A(82) and B(78)) xor (A(83) and B(77)) xor (A(84) and B(76)) xor (A(85) and B(75)) xor (A(86) and B(74)) xor (A(87) and B(73)) xor (A(88) and B(72)) xor (A(89) and B(71)) xor (A(90) and B(70)) xor (A(91) and B(69)) xor (A(92) and B(68)) xor (A(93) and B(67)) xor (A(94) and B(66)) xor (A(95) and B(65)) xor (A(96) and B(64)) xor (A(97) and B(63)) xor (A(98) and B(62)) xor (A(99) and B(61)) xor (A(100) and B(60)) xor (A(101) and B(59)) xor (A(102) and B(58)) xor (A(103) and B(57)) xor (A(104) and B(56)) xor (A(105) and B(55)) xor (A(106) and B(54)) xor (A(107) and B(53)) xor (A(108) and B(52)) xor (A(109) and B(51)) xor (A(110) and B(50)) xor (A(111) and B(49)) xor (A(112) and B(48)) xor (A(113) and B(47)) xor (A(114) and B(46)) xor (A(115) and B(45)) xor (A(116) and B(44)) xor (A(117) and B(43)) xor (A(118) and B(42)) xor (A(119) and B(41)) xor (A(120) and B(40)) xor (A(121) and B(39)) xor (A(122) and B(38)) xor (A(123) and B(37)) xor (A(124) and B(36)) xor (A(125) and B(35)) xor (A(126) and B(35));
    C(34)  <= (A(0) and B(34)) xor (A(1) and B(33)) xor (A(2) and B(32)) xor (A(3) and B(31)) xor (A(4) and B(30)) xor (A(5) and B(29)) xor (A(6) and B(28)) xor (A(7) and B(27)) xor (A(8) and B(26)) xor (A(9) and B(25)) xor (A(10) and B(24)) xor (A(11) and B(23)) xor (A(12) and B(23)) xor (A(13) and B(21)) xor (A(14) and B(20)) xor (A(15) and B(19)) xor (A(16) and B(18)) xor (A(17) and B(17)) xor (A(18) and B(16)) xor (A(19) and B(15)) xor (A(20) and B(14)) xor (A(21) and B(13)) xor (A(23) and B(12)) xor (A(23) and B(11)) xor (A(24) and B(10)) xor (A(25) and B(9)) xor (A(26) and B(8)) xor (A(27) and B(7)) xor (A(28) and B(6)) xor (A(29) and B(5)) xor (A(30) and B(4)) xor (A(31) and B(3)) xor (A(32) and B(2)) xor (A(33) and B(1)) xor (A(34) and B(0)) xor (A(27) and B(127)) xor (A(28) and B(126)) xor (A(29) and B(125)) xor (A(30) and B(124)) xor (A(31) and B(123)) xor (A(32) and B(122)) xor (A(33) and B(121)) xor (A(34) and B(120)) xor (A(35) and B(119)) xor (A(36) and B(118)) xor (A(37) and B(117)) xor (A(38) and B(116)) xor (A(39) and B(115)) xor (A(40) and B(114)) xor (A(41) and B(113)) xor (A(42) and B(112)) xor (A(43) and B(111)) xor (A(44) and B(110)) xor (A(45) and B(109)) xor (A(46) and B(108)) xor (A(47) and B(107)) xor (A(48) and B(106)) xor (A(49) and B(105)) xor (A(50) and B(104)) xor (A(51) and B(103)) xor (A(52) and B(102)) xor (A(53) and B(101)) xor (A(54) and B(100)) xor (A(55) and B(99)) xor (A(56) and B(98)) xor (A(57) and B(97)) xor (A(58) and B(96)) xor (A(59) and B(95)) xor (A(60) and B(94)) xor (A(61) and B(93)) xor (A(62) and B(92)) xor (A(63) and B(91)) xor (A(64) and B(90)) xor (A(65) and B(89)) xor (A(66) and B(88)) xor (A(67) and B(87)) xor (A(68) and B(86)) xor (A(69) and B(85)) xor (A(70) and B(84)) xor (A(71) and B(83)) xor (A(72) and B(82)) xor (A(73) and B(81)) xor (A(74) and B(80)) xor (A(75) and B(79)) xor (A(76) and B(78)) xor (A(77) and B(77)) xor (A(78) and B(76)) xor (A(79) and B(75)) xor (A(80) and B(74)) xor (A(81) and B(73)) xor (A(82) and B(72)) xor (A(83) and B(71)) xor (A(84) and B(70)) xor (A(85) and B(69)) xor (A(86) and B(68)) xor (A(87) and B(67)) xor (A(88) and B(66)) xor (A(89) and B(65)) xor (A(90) and B(64)) xor (A(91) and B(63)) xor (A(92) and B(62)) xor (A(93) and B(61)) xor (A(94) and B(60)) xor (A(95) and B(59)) xor (A(96) and B(58)) xor (A(97) and B(57)) xor (A(98) and B(56)) xor (A(99) and B(55)) xor (A(100) and B(54)) xor (A(101) and B(53)) xor (A(102) and B(52)) xor (A(103) and B(51)) xor (A(104) and B(50)) xor (A(105) and B(49)) xor (A(106) and B(48)) xor (A(107) and B(47)) xor (A(108) and B(46)) xor (A(109) and B(45)) xor (A(110) and B(44)) xor (A(111) and B(43)) xor (A(112) and B(42)) xor (A(113) and B(41)) xor (A(114) and B(40)) xor (A(115) and B(39)) xor (A(116) and B(38)) xor (A(117) and B(37)) xor (A(118) and B(36)) xor (A(119) and B(35)) xor (A(120) and B(34)) xor (A(121) and B(33)) xor (A(122) and B(32)) xor (A(123) and B(31)) xor (A(124) and B(30)) xor (A(125) and B(29)) xor (A(126) and B(28)) xor (A(32) and B(127)) xor (A(33) and B(126)) xor (A(34) and B(125)) xor (A(35) and B(124)) xor (A(36) and B(123)) xor (A(37) and B(122)) xor (A(38) and B(121)) xor (A(39) and B(120)) xor (A(40) and B(119)) xor (A(41) and B(118)) xor (A(42) and B(117)) xor (A(43) and B(116)) xor (A(44) and B(115)) xor (A(45) and B(114)) xor (A(46) and B(113)) xor (A(47) and B(112)) xor (A(48) and B(111)) xor (A(49) and B(110)) xor (A(50) and B(109)) xor (A(51) and B(108)) xor (A(52) and B(107)) xor (A(53) and B(106)) xor (A(54) and B(105)) xor (A(55) and B(104)) xor (A(56) and B(103)) xor (A(57) and B(102)) xor (A(58) and B(101)) xor (A(59) and B(100)) xor (A(60) and B(99)) xor (A(61) and B(98)) xor (A(62) and B(97)) xor (A(63) and B(96)) xor (A(64) and B(95)) xor (A(65) and B(94)) xor (A(66) and B(93)) xor (A(67) and B(92)) xor (A(68) and B(91)) xor (A(69) and B(90)) xor (A(70) and B(89)) xor (A(71) and B(88)) xor (A(72) and B(87)) xor (A(73) and B(86)) xor (A(74) and B(85)) xor (A(75) and B(84)) xor (A(76) and B(83)) xor (A(77) and B(82)) xor (A(78) and B(81)) xor (A(79) and B(80)) xor (A(80) and B(79)) xor (A(81) and B(78)) xor (A(82) and B(77)) xor (A(83) and B(76)) xor (A(84) and B(75)) xor (A(85) and B(74)) xor (A(86) and B(73)) xor (A(87) and B(72)) xor (A(88) and B(71)) xor (A(89) and B(70)) xor (A(90) and B(69)) xor (A(91) and B(68)) xor (A(92) and B(67)) xor (A(93) and B(66)) xor (A(94) and B(65)) xor (A(95) and B(64)) xor (A(96) and B(63)) xor (A(97) and B(62)) xor (A(98) and B(61)) xor (A(99) and B(60)) xor (A(100) and B(59)) xor (A(101) and B(58)) xor (A(102) and B(57)) xor (A(103) and B(56)) xor (A(104) and B(55)) xor (A(105) and B(54)) xor (A(106) and B(53)) xor (A(107) and B(52)) xor (A(108) and B(51)) xor (A(109) and B(50)) xor (A(110) and B(49)) xor (A(111) and B(48)) xor (A(112) and B(47)) xor (A(113) and B(46)) xor (A(114) and B(45)) xor (A(115) and B(44)) xor (A(116) and B(43)) xor (A(117) and B(42)) xor (A(118) and B(41)) xor (A(119) and B(40)) xor (A(120) and B(39)) xor (A(121) and B(38)) xor (A(122) and B(37)) xor (A(123) and B(36)) xor (A(124) and B(35)) xor (A(125) and B(34)) xor (A(126) and B(33)) xor (A(33) and B(127)) xor (A(34) and B(126)) xor (A(35) and B(125)) xor (A(36) and B(124)) xor (A(37) and B(123)) xor (A(38) and B(122)) xor (A(39) and B(121)) xor (A(40) and B(120)) xor (A(41) and B(119)) xor (A(42) and B(118)) xor (A(43) and B(117)) xor (A(44) and B(116)) xor (A(45) and B(115)) xor (A(46) and B(114)) xor (A(47) and B(113)) xor (A(48) and B(112)) xor (A(49) and B(111)) xor (A(50) and B(110)) xor (A(51) and B(109)) xor (A(52) and B(108)) xor (A(53) and B(107)) xor (A(54) and B(106)) xor (A(55) and B(105)) xor (A(56) and B(104)) xor (A(57) and B(103)) xor (A(58) and B(102)) xor (A(59) and B(101)) xor (A(60) and B(100)) xor (A(61) and B(99)) xor (A(62) and B(98)) xor (A(63) and B(97)) xor (A(64) and B(96)) xor (A(65) and B(95)) xor (A(66) and B(94)) xor (A(67) and B(93)) xor (A(68) and B(92)) xor (A(69) and B(91)) xor (A(70) and B(90)) xor (A(71) and B(89)) xor (A(72) and B(88)) xor (A(73) and B(87)) xor (A(74) and B(86)) xor (A(75) and B(85)) xor (A(76) and B(84)) xor (A(77) and B(83)) xor (A(78) and B(82)) xor (A(79) and B(81)) xor (A(80) and B(80)) xor (A(81) and B(79)) xor (A(82) and B(78)) xor (A(83) and B(77)) xor (A(84) and B(76)) xor (A(85) and B(75)) xor (A(86) and B(74)) xor (A(87) and B(73)) xor (A(88) and B(72)) xor (A(89) and B(71)) xor (A(90) and B(70)) xor (A(91) and B(69)) xor (A(92) and B(68)) xor (A(93) and B(67)) xor (A(94) and B(66)) xor (A(95) and B(65)) xor (A(96) and B(64)) xor (A(97) and B(63)) xor (A(98) and B(62)) xor (A(99) and B(61)) xor (A(100) and B(60)) xor (A(101) and B(59)) xor (A(102) and B(58)) xor (A(103) and B(57)) xor (A(104) and B(56)) xor (A(105) and B(55)) xor (A(106) and B(54)) xor (A(107) and B(53)) xor (A(108) and B(52)) xor (A(109) and B(51)) xor (A(110) and B(50)) xor (A(111) and B(49)) xor (A(112) and B(48)) xor (A(113) and B(47)) xor (A(114) and B(46)) xor (A(115) and B(45)) xor (A(116) and B(44)) xor (A(117) and B(43)) xor (A(118) and B(42)) xor (A(119) and B(41)) xor (A(120) and B(40)) xor (A(121) and B(39)) xor (A(122) and B(38)) xor (A(123) and B(37)) xor (A(124) and B(36)) xor (A(125) and B(35)) xor (A(126) and B(34)) xor (A(34) and B(127)) xor (A(35) and B(126)) xor (A(36) and B(125)) xor (A(37) and B(124)) xor (A(38) and B(123)) xor (A(39) and B(122)) xor (A(40) and B(121)) xor (A(41) and B(120)) xor (A(42) and B(119)) xor (A(43) and B(118)) xor (A(44) and B(117)) xor (A(45) and B(116)) xor (A(46) and B(115)) xor (A(47) and B(114)) xor (A(48) and B(113)) xor (A(49) and B(112)) xor (A(50) and B(111)) xor (A(51) and B(110)) xor (A(52) and B(109)) xor (A(53) and B(108)) xor (A(54) and B(107)) xor (A(55) and B(106)) xor (A(56) and B(105)) xor (A(57) and B(104)) xor (A(58) and B(103)) xor (A(59) and B(102)) xor (A(60) and B(101)) xor (A(61) and B(100)) xor (A(62) and B(99)) xor (A(63) and B(98)) xor (A(64) and B(97)) xor (A(65) and B(96)) xor (A(66) and B(95)) xor (A(67) and B(94)) xor (A(68) and B(93)) xor (A(69) and B(92)) xor (A(70) and B(91)) xor (A(71) and B(90)) xor (A(72) and B(89)) xor (A(73) and B(88)) xor (A(74) and B(87)) xor (A(75) and B(86)) xor (A(76) and B(85)) xor (A(77) and B(84)) xor (A(78) and B(83)) xor (A(79) and B(82)) xor (A(80) and B(81)) xor (A(81) and B(80)) xor (A(82) and B(79)) xor (A(83) and B(78)) xor (A(84) and B(77)) xor (A(85) and B(76)) xor (A(86) and B(75)) xor (A(87) and B(74)) xor (A(88) and B(73)) xor (A(89) and B(72)) xor (A(90) and B(71)) xor (A(91) and B(70)) xor (A(92) and B(69)) xor (A(93) and B(68)) xor (A(94) and B(67)) xor (A(95) and B(66)) xor (A(96) and B(65)) xor (A(97) and B(64)) xor (A(98) and B(63)) xor (A(99) and B(62)) xor (A(100) and B(61)) xor (A(101) and B(60)) xor (A(102) and B(59)) xor (A(103) and B(58)) xor (A(104) and B(57)) xor (A(105) and B(56)) xor (A(106) and B(55)) xor (A(107) and B(54)) xor (A(108) and B(53)) xor (A(109) and B(52)) xor (A(110) and B(51)) xor (A(111) and B(50)) xor (A(112) and B(49)) xor (A(113) and B(48)) xor (A(114) and B(47)) xor (A(115) and B(46)) xor (A(116) and B(45)) xor (A(117) and B(44)) xor (A(118) and B(43)) xor (A(119) and B(42)) xor (A(120) and B(41)) xor (A(121) and B(40)) xor (A(122) and B(39)) xor (A(123) and B(38)) xor (A(124) and B(37)) xor (A(125) and B(36)) xor (A(126) and B(36));
    C(35)  <= (A(0) and B(35)) xor (A(1) and B(34)) xor (A(2) and B(33)) xor (A(3) and B(32)) xor (A(4) and B(31)) xor (A(5) and B(30)) xor (A(6) and B(29)) xor (A(7) and B(28)) xor (A(8) and B(27)) xor (A(9) and B(26)) xor (A(10) and B(25)) xor (A(11) and B(24)) xor (A(12) and B(23)) xor (A(13) and B(23)) xor (A(14) and B(21)) xor (A(15) and B(20)) xor (A(16) and B(19)) xor (A(17) and B(18)) xor (A(18) and B(17)) xor (A(19) and B(16)) xor (A(20) and B(15)) xor (A(21) and B(14)) xor (A(23) and B(13)) xor (A(23) and B(12)) xor (A(24) and B(11)) xor (A(25) and B(10)) xor (A(26) and B(9)) xor (A(27) and B(8)) xor (A(28) and B(7)) xor (A(29) and B(6)) xor (A(30) and B(5)) xor (A(31) and B(4)) xor (A(32) and B(3)) xor (A(33) and B(2)) xor (A(34) and B(1)) xor (A(35) and B(0)) xor (A(28) and B(127)) xor (A(29) and B(126)) xor (A(30) and B(125)) xor (A(31) and B(124)) xor (A(32) and B(123)) xor (A(33) and B(122)) xor (A(34) and B(121)) xor (A(35) and B(120)) xor (A(36) and B(119)) xor (A(37) and B(118)) xor (A(38) and B(117)) xor (A(39) and B(116)) xor (A(40) and B(115)) xor (A(41) and B(114)) xor (A(42) and B(113)) xor (A(43) and B(112)) xor (A(44) and B(111)) xor (A(45) and B(110)) xor (A(46) and B(109)) xor (A(47) and B(108)) xor (A(48) and B(107)) xor (A(49) and B(106)) xor (A(50) and B(105)) xor (A(51) and B(104)) xor (A(52) and B(103)) xor (A(53) and B(102)) xor (A(54) and B(101)) xor (A(55) and B(100)) xor (A(56) and B(99)) xor (A(57) and B(98)) xor (A(58) and B(97)) xor (A(59) and B(96)) xor (A(60) and B(95)) xor (A(61) and B(94)) xor (A(62) and B(93)) xor (A(63) and B(92)) xor (A(64) and B(91)) xor (A(65) and B(90)) xor (A(66) and B(89)) xor (A(67) and B(88)) xor (A(68) and B(87)) xor (A(69) and B(86)) xor (A(70) and B(85)) xor (A(71) and B(84)) xor (A(72) and B(83)) xor (A(73) and B(82)) xor (A(74) and B(81)) xor (A(75) and B(80)) xor (A(76) and B(79)) xor (A(77) and B(78)) xor (A(78) and B(77)) xor (A(79) and B(76)) xor (A(80) and B(75)) xor (A(81) and B(74)) xor (A(82) and B(73)) xor (A(83) and B(72)) xor (A(84) and B(71)) xor (A(85) and B(70)) xor (A(86) and B(69)) xor (A(87) and B(68)) xor (A(88) and B(67)) xor (A(89) and B(66)) xor (A(90) and B(65)) xor (A(91) and B(64)) xor (A(92) and B(63)) xor (A(93) and B(62)) xor (A(94) and B(61)) xor (A(95) and B(60)) xor (A(96) and B(59)) xor (A(97) and B(58)) xor (A(98) and B(57)) xor (A(99) and B(56)) xor (A(100) and B(55)) xor (A(101) and B(54)) xor (A(102) and B(53)) xor (A(103) and B(52)) xor (A(104) and B(51)) xor (A(105) and B(50)) xor (A(106) and B(49)) xor (A(107) and B(48)) xor (A(108) and B(47)) xor (A(109) and B(46)) xor (A(110) and B(45)) xor (A(111) and B(44)) xor (A(112) and B(43)) xor (A(113) and B(42)) xor (A(114) and B(41)) xor (A(115) and B(40)) xor (A(116) and B(39)) xor (A(117) and B(38)) xor (A(118) and B(37)) xor (A(119) and B(36)) xor (A(120) and B(35)) xor (A(121) and B(34)) xor (A(122) and B(33)) xor (A(123) and B(32)) xor (A(124) and B(31)) xor (A(125) and B(30)) xor (A(126) and B(29)) xor (A(33) and B(127)) xor (A(34) and B(126)) xor (A(35) and B(125)) xor (A(36) and B(124)) xor (A(37) and B(123)) xor (A(38) and B(122)) xor (A(39) and B(121)) xor (A(40) and B(120)) xor (A(41) and B(119)) xor (A(42) and B(118)) xor (A(43) and B(117)) xor (A(44) and B(116)) xor (A(45) and B(115)) xor (A(46) and B(114)) xor (A(47) and B(113)) xor (A(48) and B(112)) xor (A(49) and B(111)) xor (A(50) and B(110)) xor (A(51) and B(109)) xor (A(52) and B(108)) xor (A(53) and B(107)) xor (A(54) and B(106)) xor (A(55) and B(105)) xor (A(56) and B(104)) xor (A(57) and B(103)) xor (A(58) and B(102)) xor (A(59) and B(101)) xor (A(60) and B(100)) xor (A(61) and B(99)) xor (A(62) and B(98)) xor (A(63) and B(97)) xor (A(64) and B(96)) xor (A(65) and B(95)) xor (A(66) and B(94)) xor (A(67) and B(93)) xor (A(68) and B(92)) xor (A(69) and B(91)) xor (A(70) and B(90)) xor (A(71) and B(89)) xor (A(72) and B(88)) xor (A(73) and B(87)) xor (A(74) and B(86)) xor (A(75) and B(85)) xor (A(76) and B(84)) xor (A(77) and B(83)) xor (A(78) and B(82)) xor (A(79) and B(81)) xor (A(80) and B(80)) xor (A(81) and B(79)) xor (A(82) and B(78)) xor (A(83) and B(77)) xor (A(84) and B(76)) xor (A(85) and B(75)) xor (A(86) and B(74)) xor (A(87) and B(73)) xor (A(88) and B(72)) xor (A(89) and B(71)) xor (A(90) and B(70)) xor (A(91) and B(69)) xor (A(92) and B(68)) xor (A(93) and B(67)) xor (A(94) and B(66)) xor (A(95) and B(65)) xor (A(96) and B(64)) xor (A(97) and B(63)) xor (A(98) and B(62)) xor (A(99) and B(61)) xor (A(100) and B(60)) xor (A(101) and B(59)) xor (A(102) and B(58)) xor (A(103) and B(57)) xor (A(104) and B(56)) xor (A(105) and B(55)) xor (A(106) and B(54)) xor (A(107) and B(53)) xor (A(108) and B(52)) xor (A(109) and B(51)) xor (A(110) and B(50)) xor (A(111) and B(49)) xor (A(112) and B(48)) xor (A(113) and B(47)) xor (A(114) and B(46)) xor (A(115) and B(45)) xor (A(116) and B(44)) xor (A(117) and B(43)) xor (A(118) and B(42)) xor (A(119) and B(41)) xor (A(120) and B(40)) xor (A(121) and B(39)) xor (A(122) and B(38)) xor (A(123) and B(37)) xor (A(124) and B(36)) xor (A(125) and B(35)) xor (A(126) and B(34)) xor (A(34) and B(127)) xor (A(35) and B(126)) xor (A(36) and B(125)) xor (A(37) and B(124)) xor (A(38) and B(123)) xor (A(39) and B(122)) xor (A(40) and B(121)) xor (A(41) and B(120)) xor (A(42) and B(119)) xor (A(43) and B(118)) xor (A(44) and B(117)) xor (A(45) and B(116)) xor (A(46) and B(115)) xor (A(47) and B(114)) xor (A(48) and B(113)) xor (A(49) and B(112)) xor (A(50) and B(111)) xor (A(51) and B(110)) xor (A(52) and B(109)) xor (A(53) and B(108)) xor (A(54) and B(107)) xor (A(55) and B(106)) xor (A(56) and B(105)) xor (A(57) and B(104)) xor (A(58) and B(103)) xor (A(59) and B(102)) xor (A(60) and B(101)) xor (A(61) and B(100)) xor (A(62) and B(99)) xor (A(63) and B(98)) xor (A(64) and B(97)) xor (A(65) and B(96)) xor (A(66) and B(95)) xor (A(67) and B(94)) xor (A(68) and B(93)) xor (A(69) and B(92)) xor (A(70) and B(91)) xor (A(71) and B(90)) xor (A(72) and B(89)) xor (A(73) and B(88)) xor (A(74) and B(87)) xor (A(75) and B(86)) xor (A(76) and B(85)) xor (A(77) and B(84)) xor (A(78) and B(83)) xor (A(79) and B(82)) xor (A(80) and B(81)) xor (A(81) and B(80)) xor (A(82) and B(79)) xor (A(83) and B(78)) xor (A(84) and B(77)) xor (A(85) and B(76)) xor (A(86) and B(75)) xor (A(87) and B(74)) xor (A(88) and B(73)) xor (A(89) and B(72)) xor (A(90) and B(71)) xor (A(91) and B(70)) xor (A(92) and B(69)) xor (A(93) and B(68)) xor (A(94) and B(67)) xor (A(95) and B(66)) xor (A(96) and B(65)) xor (A(97) and B(64)) xor (A(98) and B(63)) xor (A(99) and B(62)) xor (A(100) and B(61)) xor (A(101) and B(60)) xor (A(102) and B(59)) xor (A(103) and B(58)) xor (A(104) and B(57)) xor (A(105) and B(56)) xor (A(106) and B(55)) xor (A(107) and B(54)) xor (A(108) and B(53)) xor (A(109) and B(52)) xor (A(110) and B(51)) xor (A(111) and B(50)) xor (A(112) and B(49)) xor (A(113) and B(48)) xor (A(114) and B(47)) xor (A(115) and B(46)) xor (A(116) and B(45)) xor (A(117) and B(44)) xor (A(118) and B(43)) xor (A(119) and B(42)) xor (A(120) and B(41)) xor (A(121) and B(40)) xor (A(122) and B(39)) xor (A(123) and B(38)) xor (A(124) and B(37)) xor (A(125) and B(36)) xor (A(126) and B(35)) xor (A(35) and B(127)) xor (A(36) and B(126)) xor (A(37) and B(125)) xor (A(38) and B(124)) xor (A(39) and B(123)) xor (A(40) and B(122)) xor (A(41) and B(121)) xor (A(42) and B(120)) xor (A(43) and B(119)) xor (A(44) and B(118)) xor (A(45) and B(117)) xor (A(46) and B(116)) xor (A(47) and B(115)) xor (A(48) and B(114)) xor (A(49) and B(113)) xor (A(50) and B(112)) xor (A(51) and B(111)) xor (A(52) and B(110)) xor (A(53) and B(109)) xor (A(54) and B(108)) xor (A(55) and B(107)) xor (A(56) and B(106)) xor (A(57) and B(105)) xor (A(58) and B(104)) xor (A(59) and B(103)) xor (A(60) and B(102)) xor (A(61) and B(101)) xor (A(62) and B(100)) xor (A(63) and B(99)) xor (A(64) and B(98)) xor (A(65) and B(97)) xor (A(66) and B(96)) xor (A(67) and B(95)) xor (A(68) and B(94)) xor (A(69) and B(93)) xor (A(70) and B(92)) xor (A(71) and B(91)) xor (A(72) and B(90)) xor (A(73) and B(89)) xor (A(74) and B(88)) xor (A(75) and B(87)) xor (A(76) and B(86)) xor (A(77) and B(85)) xor (A(78) and B(84)) xor (A(79) and B(83)) xor (A(80) and B(82)) xor (A(81) and B(81)) xor (A(82) and B(80)) xor (A(83) and B(79)) xor (A(84) and B(78)) xor (A(85) and B(77)) xor (A(86) and B(76)) xor (A(87) and B(75)) xor (A(88) and B(74)) xor (A(89) and B(73)) xor (A(90) and B(72)) xor (A(91) and B(71)) xor (A(92) and B(70)) xor (A(93) and B(69)) xor (A(94) and B(68)) xor (A(95) and B(67)) xor (A(96) and B(66)) xor (A(97) and B(65)) xor (A(98) and B(64)) xor (A(99) and B(63)) xor (A(100) and B(62)) xor (A(101) and B(61)) xor (A(102) and B(60)) xor (A(103) and B(59)) xor (A(104) and B(58)) xor (A(105) and B(57)) xor (A(106) and B(56)) xor (A(107) and B(55)) xor (A(108) and B(54)) xor (A(109) and B(53)) xor (A(110) and B(52)) xor (A(111) and B(51)) xor (A(112) and B(50)) xor (A(113) and B(49)) xor (A(114) and B(48)) xor (A(115) and B(47)) xor (A(116) and B(46)) xor (A(117) and B(45)) xor (A(118) and B(44)) xor (A(119) and B(43)) xor (A(120) and B(42)) xor (A(121) and B(41)) xor (A(122) and B(40)) xor (A(123) and B(39)) xor (A(124) and B(38)) xor (A(125) and B(37)) xor (A(126) and B(37));
    C(36)  <= (A(0) and B(36)) xor (A(1) and B(35)) xor (A(2) and B(34)) xor (A(3) and B(33)) xor (A(4) and B(32)) xor (A(5) and B(31)) xor (A(6) and B(30)) xor (A(7) and B(29)) xor (A(8) and B(28)) xor (A(9) and B(27)) xor (A(10) and B(26)) xor (A(11) and B(25)) xor (A(12) and B(24)) xor (A(13) and B(23)) xor (A(14) and B(23)) xor (A(15) and B(21)) xor (A(16) and B(20)) xor (A(17) and B(19)) xor (A(18) and B(18)) xor (A(19) and B(17)) xor (A(20) and B(16)) xor (A(21) and B(15)) xor (A(23) and B(14)) xor (A(23) and B(13)) xor (A(24) and B(12)) xor (A(25) and B(11)) xor (A(26) and B(10)) xor (A(27) and B(9)) xor (A(28) and B(8)) xor (A(29) and B(7)) xor (A(30) and B(6)) xor (A(31) and B(5)) xor (A(32) and B(4)) xor (A(33) and B(3)) xor (A(34) and B(2)) xor (A(35) and B(1)) xor (A(36) and B(0)) xor (A(29) and B(127)) xor (A(30) and B(126)) xor (A(31) and B(125)) xor (A(32) and B(124)) xor (A(33) and B(123)) xor (A(34) and B(122)) xor (A(35) and B(121)) xor (A(36) and B(120)) xor (A(37) and B(119)) xor (A(38) and B(118)) xor (A(39) and B(117)) xor (A(40) and B(116)) xor (A(41) and B(115)) xor (A(42) and B(114)) xor (A(43) and B(113)) xor (A(44) and B(112)) xor (A(45) and B(111)) xor (A(46) and B(110)) xor (A(47) and B(109)) xor (A(48) and B(108)) xor (A(49) and B(107)) xor (A(50) and B(106)) xor (A(51) and B(105)) xor (A(52) and B(104)) xor (A(53) and B(103)) xor (A(54) and B(102)) xor (A(55) and B(101)) xor (A(56) and B(100)) xor (A(57) and B(99)) xor (A(58) and B(98)) xor (A(59) and B(97)) xor (A(60) and B(96)) xor (A(61) and B(95)) xor (A(62) and B(94)) xor (A(63) and B(93)) xor (A(64) and B(92)) xor (A(65) and B(91)) xor (A(66) and B(90)) xor (A(67) and B(89)) xor (A(68) and B(88)) xor (A(69) and B(87)) xor (A(70) and B(86)) xor (A(71) and B(85)) xor (A(72) and B(84)) xor (A(73) and B(83)) xor (A(74) and B(82)) xor (A(75) and B(81)) xor (A(76) and B(80)) xor (A(77) and B(79)) xor (A(78) and B(78)) xor (A(79) and B(77)) xor (A(80) and B(76)) xor (A(81) and B(75)) xor (A(82) and B(74)) xor (A(83) and B(73)) xor (A(84) and B(72)) xor (A(85) and B(71)) xor (A(86) and B(70)) xor (A(87) and B(69)) xor (A(88) and B(68)) xor (A(89) and B(67)) xor (A(90) and B(66)) xor (A(91) and B(65)) xor (A(92) and B(64)) xor (A(93) and B(63)) xor (A(94) and B(62)) xor (A(95) and B(61)) xor (A(96) and B(60)) xor (A(97) and B(59)) xor (A(98) and B(58)) xor (A(99) and B(57)) xor (A(100) and B(56)) xor (A(101) and B(55)) xor (A(102) and B(54)) xor (A(103) and B(53)) xor (A(104) and B(52)) xor (A(105) and B(51)) xor (A(106) and B(50)) xor (A(107) and B(49)) xor (A(108) and B(48)) xor (A(109) and B(47)) xor (A(110) and B(46)) xor (A(111) and B(45)) xor (A(112) and B(44)) xor (A(113) and B(43)) xor (A(114) and B(42)) xor (A(115) and B(41)) xor (A(116) and B(40)) xor (A(117) and B(39)) xor (A(118) and B(38)) xor (A(119) and B(37)) xor (A(120) and B(36)) xor (A(121) and B(35)) xor (A(122) and B(34)) xor (A(123) and B(33)) xor (A(124) and B(32)) xor (A(125) and B(31)) xor (A(126) and B(30)) xor (A(34) and B(127)) xor (A(35) and B(126)) xor (A(36) and B(125)) xor (A(37) and B(124)) xor (A(38) and B(123)) xor (A(39) and B(122)) xor (A(40) and B(121)) xor (A(41) and B(120)) xor (A(42) and B(119)) xor (A(43) and B(118)) xor (A(44) and B(117)) xor (A(45) and B(116)) xor (A(46) and B(115)) xor (A(47) and B(114)) xor (A(48) and B(113)) xor (A(49) and B(112)) xor (A(50) and B(111)) xor (A(51) and B(110)) xor (A(52) and B(109)) xor (A(53) and B(108)) xor (A(54) and B(107)) xor (A(55) and B(106)) xor (A(56) and B(105)) xor (A(57) and B(104)) xor (A(58) and B(103)) xor (A(59) and B(102)) xor (A(60) and B(101)) xor (A(61) and B(100)) xor (A(62) and B(99)) xor (A(63) and B(98)) xor (A(64) and B(97)) xor (A(65) and B(96)) xor (A(66) and B(95)) xor (A(67) and B(94)) xor (A(68) and B(93)) xor (A(69) and B(92)) xor (A(70) and B(91)) xor (A(71) and B(90)) xor (A(72) and B(89)) xor (A(73) and B(88)) xor (A(74) and B(87)) xor (A(75) and B(86)) xor (A(76) and B(85)) xor (A(77) and B(84)) xor (A(78) and B(83)) xor (A(79) and B(82)) xor (A(80) and B(81)) xor (A(81) and B(80)) xor (A(82) and B(79)) xor (A(83) and B(78)) xor (A(84) and B(77)) xor (A(85) and B(76)) xor (A(86) and B(75)) xor (A(87) and B(74)) xor (A(88) and B(73)) xor (A(89) and B(72)) xor (A(90) and B(71)) xor (A(91) and B(70)) xor (A(92) and B(69)) xor (A(93) and B(68)) xor (A(94) and B(67)) xor (A(95) and B(66)) xor (A(96) and B(65)) xor (A(97) and B(64)) xor (A(98) and B(63)) xor (A(99) and B(62)) xor (A(100) and B(61)) xor (A(101) and B(60)) xor (A(102) and B(59)) xor (A(103) and B(58)) xor (A(104) and B(57)) xor (A(105) and B(56)) xor (A(106) and B(55)) xor (A(107) and B(54)) xor (A(108) and B(53)) xor (A(109) and B(52)) xor (A(110) and B(51)) xor (A(111) and B(50)) xor (A(112) and B(49)) xor (A(113) and B(48)) xor (A(114) and B(47)) xor (A(115) and B(46)) xor (A(116) and B(45)) xor (A(117) and B(44)) xor (A(118) and B(43)) xor (A(119) and B(42)) xor (A(120) and B(41)) xor (A(121) and B(40)) xor (A(122) and B(39)) xor (A(123) and B(38)) xor (A(124) and B(37)) xor (A(125) and B(36)) xor (A(126) and B(35)) xor (A(35) and B(127)) xor (A(36) and B(126)) xor (A(37) and B(125)) xor (A(38) and B(124)) xor (A(39) and B(123)) xor (A(40) and B(122)) xor (A(41) and B(121)) xor (A(42) and B(120)) xor (A(43) and B(119)) xor (A(44) and B(118)) xor (A(45) and B(117)) xor (A(46) and B(116)) xor (A(47) and B(115)) xor (A(48) and B(114)) xor (A(49) and B(113)) xor (A(50) and B(112)) xor (A(51) and B(111)) xor (A(52) and B(110)) xor (A(53) and B(109)) xor (A(54) and B(108)) xor (A(55) and B(107)) xor (A(56) and B(106)) xor (A(57) and B(105)) xor (A(58) and B(104)) xor (A(59) and B(103)) xor (A(60) and B(102)) xor (A(61) and B(101)) xor (A(62) and B(100)) xor (A(63) and B(99)) xor (A(64) and B(98)) xor (A(65) and B(97)) xor (A(66) and B(96)) xor (A(67) and B(95)) xor (A(68) and B(94)) xor (A(69) and B(93)) xor (A(70) and B(92)) xor (A(71) and B(91)) xor (A(72) and B(90)) xor (A(73) and B(89)) xor (A(74) and B(88)) xor (A(75) and B(87)) xor (A(76) and B(86)) xor (A(77) and B(85)) xor (A(78) and B(84)) xor (A(79) and B(83)) xor (A(80) and B(82)) xor (A(81) and B(81)) xor (A(82) and B(80)) xor (A(83) and B(79)) xor (A(84) and B(78)) xor (A(85) and B(77)) xor (A(86) and B(76)) xor (A(87) and B(75)) xor (A(88) and B(74)) xor (A(89) and B(73)) xor (A(90) and B(72)) xor (A(91) and B(71)) xor (A(92) and B(70)) xor (A(93) and B(69)) xor (A(94) and B(68)) xor (A(95) and B(67)) xor (A(96) and B(66)) xor (A(97) and B(65)) xor (A(98) and B(64)) xor (A(99) and B(63)) xor (A(100) and B(62)) xor (A(101) and B(61)) xor (A(102) and B(60)) xor (A(103) and B(59)) xor (A(104) and B(58)) xor (A(105) and B(57)) xor (A(106) and B(56)) xor (A(107) and B(55)) xor (A(108) and B(54)) xor (A(109) and B(53)) xor (A(110) and B(52)) xor (A(111) and B(51)) xor (A(112) and B(50)) xor (A(113) and B(49)) xor (A(114) and B(48)) xor (A(115) and B(47)) xor (A(116) and B(46)) xor (A(117) and B(45)) xor (A(118) and B(44)) xor (A(119) and B(43)) xor (A(120) and B(42)) xor (A(121) and B(41)) xor (A(122) and B(40)) xor (A(123) and B(39)) xor (A(124) and B(38)) xor (A(125) and B(37)) xor (A(126) and B(36)) xor (A(36) and B(127)) xor (A(37) and B(126)) xor (A(38) and B(125)) xor (A(39) and B(124)) xor (A(40) and B(123)) xor (A(41) and B(122)) xor (A(42) and B(121)) xor (A(43) and B(120)) xor (A(44) and B(119)) xor (A(45) and B(118)) xor (A(46) and B(117)) xor (A(47) and B(116)) xor (A(48) and B(115)) xor (A(49) and B(114)) xor (A(50) and B(113)) xor (A(51) and B(112)) xor (A(52) and B(111)) xor (A(53) and B(110)) xor (A(54) and B(109)) xor (A(55) and B(108)) xor (A(56) and B(107)) xor (A(57) and B(106)) xor (A(58) and B(105)) xor (A(59) and B(104)) xor (A(60) and B(103)) xor (A(61) and B(102)) xor (A(62) and B(101)) xor (A(63) and B(100)) xor (A(64) and B(99)) xor (A(65) and B(98)) xor (A(66) and B(97)) xor (A(67) and B(96)) xor (A(68) and B(95)) xor (A(69) and B(94)) xor (A(70) and B(93)) xor (A(71) and B(92)) xor (A(72) and B(91)) xor (A(73) and B(90)) xor (A(74) and B(89)) xor (A(75) and B(88)) xor (A(76) and B(87)) xor (A(77) and B(86)) xor (A(78) and B(85)) xor (A(79) and B(84)) xor (A(80) and B(83)) xor (A(81) and B(82)) xor (A(82) and B(81)) xor (A(83) and B(80)) xor (A(84) and B(79)) xor (A(85) and B(78)) xor (A(86) and B(77)) xor (A(87) and B(76)) xor (A(88) and B(75)) xor (A(89) and B(74)) xor (A(90) and B(73)) xor (A(91) and B(72)) xor (A(92) and B(71)) xor (A(93) and B(70)) xor (A(94) and B(69)) xor (A(95) and B(68)) xor (A(96) and B(67)) xor (A(97) and B(66)) xor (A(98) and B(65)) xor (A(99) and B(64)) xor (A(100) and B(63)) xor (A(101) and B(62)) xor (A(102) and B(61)) xor (A(103) and B(60)) xor (A(104) and B(59)) xor (A(105) and B(58)) xor (A(106) and B(57)) xor (A(107) and B(56)) xor (A(108) and B(55)) xor (A(109) and B(54)) xor (A(110) and B(53)) xor (A(111) and B(52)) xor (A(112) and B(51)) xor (A(113) and B(50)) xor (A(114) and B(49)) xor (A(115) and B(48)) xor (A(116) and B(47)) xor (A(117) and B(46)) xor (A(118) and B(45)) xor (A(119) and B(44)) xor (A(120) and B(43)) xor (A(121) and B(42)) xor (A(122) and B(41)) xor (A(123) and B(40)) xor (A(124) and B(39)) xor (A(125) and B(38)) xor (A(126) and B(38));
    C(37)  <= (A(0) and B(37)) xor (A(1) and B(36)) xor (A(2) and B(35)) xor (A(3) and B(34)) xor (A(4) and B(33)) xor (A(5) and B(32)) xor (A(6) and B(31)) xor (A(7) and B(30)) xor (A(8) and B(29)) xor (A(9) and B(28)) xor (A(10) and B(27)) xor (A(11) and B(26)) xor (A(12) and B(25)) xor (A(13) and B(24)) xor (A(14) and B(23)) xor (A(15) and B(23)) xor (A(16) and B(21)) xor (A(17) and B(20)) xor (A(18) and B(19)) xor (A(19) and B(18)) xor (A(20) and B(17)) xor (A(21) and B(16)) xor (A(23) and B(15)) xor (A(23) and B(14)) xor (A(24) and B(13)) xor (A(25) and B(12)) xor (A(26) and B(11)) xor (A(27) and B(10)) xor (A(28) and B(9)) xor (A(29) and B(8)) xor (A(30) and B(7)) xor (A(31) and B(6)) xor (A(32) and B(5)) xor (A(33) and B(4)) xor (A(34) and B(3)) xor (A(35) and B(2)) xor (A(36) and B(1)) xor (A(37) and B(0)) xor (A(30) and B(127)) xor (A(31) and B(126)) xor (A(32) and B(125)) xor (A(33) and B(124)) xor (A(34) and B(123)) xor (A(35) and B(122)) xor (A(36) and B(121)) xor (A(37) and B(120)) xor (A(38) and B(119)) xor (A(39) and B(118)) xor (A(40) and B(117)) xor (A(41) and B(116)) xor (A(42) and B(115)) xor (A(43) and B(114)) xor (A(44) and B(113)) xor (A(45) and B(112)) xor (A(46) and B(111)) xor (A(47) and B(110)) xor (A(48) and B(109)) xor (A(49) and B(108)) xor (A(50) and B(107)) xor (A(51) and B(106)) xor (A(52) and B(105)) xor (A(53) and B(104)) xor (A(54) and B(103)) xor (A(55) and B(102)) xor (A(56) and B(101)) xor (A(57) and B(100)) xor (A(58) and B(99)) xor (A(59) and B(98)) xor (A(60) and B(97)) xor (A(61) and B(96)) xor (A(62) and B(95)) xor (A(63) and B(94)) xor (A(64) and B(93)) xor (A(65) and B(92)) xor (A(66) and B(91)) xor (A(67) and B(90)) xor (A(68) and B(89)) xor (A(69) and B(88)) xor (A(70) and B(87)) xor (A(71) and B(86)) xor (A(72) and B(85)) xor (A(73) and B(84)) xor (A(74) and B(83)) xor (A(75) and B(82)) xor (A(76) and B(81)) xor (A(77) and B(80)) xor (A(78) and B(79)) xor (A(79) and B(78)) xor (A(80) and B(77)) xor (A(81) and B(76)) xor (A(82) and B(75)) xor (A(83) and B(74)) xor (A(84) and B(73)) xor (A(85) and B(72)) xor (A(86) and B(71)) xor (A(87) and B(70)) xor (A(88) and B(69)) xor (A(89) and B(68)) xor (A(90) and B(67)) xor (A(91) and B(66)) xor (A(92) and B(65)) xor (A(93) and B(64)) xor (A(94) and B(63)) xor (A(95) and B(62)) xor (A(96) and B(61)) xor (A(97) and B(60)) xor (A(98) and B(59)) xor (A(99) and B(58)) xor (A(100) and B(57)) xor (A(101) and B(56)) xor (A(102) and B(55)) xor (A(103) and B(54)) xor (A(104) and B(53)) xor (A(105) and B(52)) xor (A(106) and B(51)) xor (A(107) and B(50)) xor (A(108) and B(49)) xor (A(109) and B(48)) xor (A(110) and B(47)) xor (A(111) and B(46)) xor (A(112) and B(45)) xor (A(113) and B(44)) xor (A(114) and B(43)) xor (A(115) and B(42)) xor (A(116) and B(41)) xor (A(117) and B(40)) xor (A(118) and B(39)) xor (A(119) and B(38)) xor (A(120) and B(37)) xor (A(121) and B(36)) xor (A(122) and B(35)) xor (A(123) and B(34)) xor (A(124) and B(33)) xor (A(125) and B(32)) xor (A(126) and B(31)) xor (A(35) and B(127)) xor (A(36) and B(126)) xor (A(37) and B(125)) xor (A(38) and B(124)) xor (A(39) and B(123)) xor (A(40) and B(122)) xor (A(41) and B(121)) xor (A(42) and B(120)) xor (A(43) and B(119)) xor (A(44) and B(118)) xor (A(45) and B(117)) xor (A(46) and B(116)) xor (A(47) and B(115)) xor (A(48) and B(114)) xor (A(49) and B(113)) xor (A(50) and B(112)) xor (A(51) and B(111)) xor (A(52) and B(110)) xor (A(53) and B(109)) xor (A(54) and B(108)) xor (A(55) and B(107)) xor (A(56) and B(106)) xor (A(57) and B(105)) xor (A(58) and B(104)) xor (A(59) and B(103)) xor (A(60) and B(102)) xor (A(61) and B(101)) xor (A(62) and B(100)) xor (A(63) and B(99)) xor (A(64) and B(98)) xor (A(65) and B(97)) xor (A(66) and B(96)) xor (A(67) and B(95)) xor (A(68) and B(94)) xor (A(69) and B(93)) xor (A(70) and B(92)) xor (A(71) and B(91)) xor (A(72) and B(90)) xor (A(73) and B(89)) xor (A(74) and B(88)) xor (A(75) and B(87)) xor (A(76) and B(86)) xor (A(77) and B(85)) xor (A(78) and B(84)) xor (A(79) and B(83)) xor (A(80) and B(82)) xor (A(81) and B(81)) xor (A(82) and B(80)) xor (A(83) and B(79)) xor (A(84) and B(78)) xor (A(85) and B(77)) xor (A(86) and B(76)) xor (A(87) and B(75)) xor (A(88) and B(74)) xor (A(89) and B(73)) xor (A(90) and B(72)) xor (A(91) and B(71)) xor (A(92) and B(70)) xor (A(93) and B(69)) xor (A(94) and B(68)) xor (A(95) and B(67)) xor (A(96) and B(66)) xor (A(97) and B(65)) xor (A(98) and B(64)) xor (A(99) and B(63)) xor (A(100) and B(62)) xor (A(101) and B(61)) xor (A(102) and B(60)) xor (A(103) and B(59)) xor (A(104) and B(58)) xor (A(105) and B(57)) xor (A(106) and B(56)) xor (A(107) and B(55)) xor (A(108) and B(54)) xor (A(109) and B(53)) xor (A(110) and B(52)) xor (A(111) and B(51)) xor (A(112) and B(50)) xor (A(113) and B(49)) xor (A(114) and B(48)) xor (A(115) and B(47)) xor (A(116) and B(46)) xor (A(117) and B(45)) xor (A(118) and B(44)) xor (A(119) and B(43)) xor (A(120) and B(42)) xor (A(121) and B(41)) xor (A(122) and B(40)) xor (A(123) and B(39)) xor (A(124) and B(38)) xor (A(125) and B(37)) xor (A(126) and B(36)) xor (A(36) and B(127)) xor (A(37) and B(126)) xor (A(38) and B(125)) xor (A(39) and B(124)) xor (A(40) and B(123)) xor (A(41) and B(122)) xor (A(42) and B(121)) xor (A(43) and B(120)) xor (A(44) and B(119)) xor (A(45) and B(118)) xor (A(46) and B(117)) xor (A(47) and B(116)) xor (A(48) and B(115)) xor (A(49) and B(114)) xor (A(50) and B(113)) xor (A(51) and B(112)) xor (A(52) and B(111)) xor (A(53) and B(110)) xor (A(54) and B(109)) xor (A(55) and B(108)) xor (A(56) and B(107)) xor (A(57) and B(106)) xor (A(58) and B(105)) xor (A(59) and B(104)) xor (A(60) and B(103)) xor (A(61) and B(102)) xor (A(62) and B(101)) xor (A(63) and B(100)) xor (A(64) and B(99)) xor (A(65) and B(98)) xor (A(66) and B(97)) xor (A(67) and B(96)) xor (A(68) and B(95)) xor (A(69) and B(94)) xor (A(70) and B(93)) xor (A(71) and B(92)) xor (A(72) and B(91)) xor (A(73) and B(90)) xor (A(74) and B(89)) xor (A(75) and B(88)) xor (A(76) and B(87)) xor (A(77) and B(86)) xor (A(78) and B(85)) xor (A(79) and B(84)) xor (A(80) and B(83)) xor (A(81) and B(82)) xor (A(82) and B(81)) xor (A(83) and B(80)) xor (A(84) and B(79)) xor (A(85) and B(78)) xor (A(86) and B(77)) xor (A(87) and B(76)) xor (A(88) and B(75)) xor (A(89) and B(74)) xor (A(90) and B(73)) xor (A(91) and B(72)) xor (A(92) and B(71)) xor (A(93) and B(70)) xor (A(94) and B(69)) xor (A(95) and B(68)) xor (A(96) and B(67)) xor (A(97) and B(66)) xor (A(98) and B(65)) xor (A(99) and B(64)) xor (A(100) and B(63)) xor (A(101) and B(62)) xor (A(102) and B(61)) xor (A(103) and B(60)) xor (A(104) and B(59)) xor (A(105) and B(58)) xor (A(106) and B(57)) xor (A(107) and B(56)) xor (A(108) and B(55)) xor (A(109) and B(54)) xor (A(110) and B(53)) xor (A(111) and B(52)) xor (A(112) and B(51)) xor (A(113) and B(50)) xor (A(114) and B(49)) xor (A(115) and B(48)) xor (A(116) and B(47)) xor (A(117) and B(46)) xor (A(118) and B(45)) xor (A(119) and B(44)) xor (A(120) and B(43)) xor (A(121) and B(42)) xor (A(122) and B(41)) xor (A(123) and B(40)) xor (A(124) and B(39)) xor (A(125) and B(38)) xor (A(126) and B(37)) xor (A(37) and B(127)) xor (A(38) and B(126)) xor (A(39) and B(125)) xor (A(40) and B(124)) xor (A(41) and B(123)) xor (A(42) and B(122)) xor (A(43) and B(121)) xor (A(44) and B(120)) xor (A(45) and B(119)) xor (A(46) and B(118)) xor (A(47) and B(117)) xor (A(48) and B(116)) xor (A(49) and B(115)) xor (A(50) and B(114)) xor (A(51) and B(113)) xor (A(52) and B(112)) xor (A(53) and B(111)) xor (A(54) and B(110)) xor (A(55) and B(109)) xor (A(56) and B(108)) xor (A(57) and B(107)) xor (A(58) and B(106)) xor (A(59) and B(105)) xor (A(60) and B(104)) xor (A(61) and B(103)) xor (A(62) and B(102)) xor (A(63) and B(101)) xor (A(64) and B(100)) xor (A(65) and B(99)) xor (A(66) and B(98)) xor (A(67) and B(97)) xor (A(68) and B(96)) xor (A(69) and B(95)) xor (A(70) and B(94)) xor (A(71) and B(93)) xor (A(72) and B(92)) xor (A(73) and B(91)) xor (A(74) and B(90)) xor (A(75) and B(89)) xor (A(76) and B(88)) xor (A(77) and B(87)) xor (A(78) and B(86)) xor (A(79) and B(85)) xor (A(80) and B(84)) xor (A(81) and B(83)) xor (A(82) and B(82)) xor (A(83) and B(81)) xor (A(84) and B(80)) xor (A(85) and B(79)) xor (A(86) and B(78)) xor (A(87) and B(77)) xor (A(88) and B(76)) xor (A(89) and B(75)) xor (A(90) and B(74)) xor (A(91) and B(73)) xor (A(92) and B(72)) xor (A(93) and B(71)) xor (A(94) and B(70)) xor (A(95) and B(69)) xor (A(96) and B(68)) xor (A(97) and B(67)) xor (A(98) and B(66)) xor (A(99) and B(65)) xor (A(100) and B(64)) xor (A(101) and B(63)) xor (A(102) and B(62)) xor (A(103) and B(61)) xor (A(104) and B(60)) xor (A(105) and B(59)) xor (A(106) and B(58)) xor (A(107) and B(57)) xor (A(108) and B(56)) xor (A(109) and B(55)) xor (A(110) and B(54)) xor (A(111) and B(53)) xor (A(112) and B(52)) xor (A(113) and B(51)) xor (A(114) and B(50)) xor (A(115) and B(49)) xor (A(116) and B(48)) xor (A(117) and B(47)) xor (A(118) and B(46)) xor (A(119) and B(45)) xor (A(120) and B(44)) xor (A(121) and B(43)) xor (A(122) and B(42)) xor (A(123) and B(41)) xor (A(124) and B(40)) xor (A(125) and B(39)) xor (A(126) and B(39));
    C(38)  <= (A(0) and B(38)) xor (A(1) and B(37)) xor (A(2) and B(36)) xor (A(3) and B(35)) xor (A(4) and B(34)) xor (A(5) and B(33)) xor (A(6) and B(32)) xor (A(7) and B(31)) xor (A(8) and B(30)) xor (A(9) and B(29)) xor (A(10) and B(28)) xor (A(11) and B(27)) xor (A(12) and B(26)) xor (A(13) and B(25)) xor (A(14) and B(24)) xor (A(15) and B(23)) xor (A(16) and B(23)) xor (A(17) and B(21)) xor (A(18) and B(20)) xor (A(19) and B(19)) xor (A(20) and B(18)) xor (A(21) and B(17)) xor (A(23) and B(16)) xor (A(23) and B(15)) xor (A(24) and B(14)) xor (A(25) and B(13)) xor (A(26) and B(12)) xor (A(27) and B(11)) xor (A(28) and B(10)) xor (A(29) and B(9)) xor (A(30) and B(8)) xor (A(31) and B(7)) xor (A(32) and B(6)) xor (A(33) and B(5)) xor (A(34) and B(4)) xor (A(35) and B(3)) xor (A(36) and B(2)) xor (A(37) and B(1)) xor (A(38) and B(0)) xor (A(31) and B(127)) xor (A(32) and B(126)) xor (A(33) and B(125)) xor (A(34) and B(124)) xor (A(35) and B(123)) xor (A(36) and B(122)) xor (A(37) and B(121)) xor (A(38) and B(120)) xor (A(39) and B(119)) xor (A(40) and B(118)) xor (A(41) and B(117)) xor (A(42) and B(116)) xor (A(43) and B(115)) xor (A(44) and B(114)) xor (A(45) and B(113)) xor (A(46) and B(112)) xor (A(47) and B(111)) xor (A(48) and B(110)) xor (A(49) and B(109)) xor (A(50) and B(108)) xor (A(51) and B(107)) xor (A(52) and B(106)) xor (A(53) and B(105)) xor (A(54) and B(104)) xor (A(55) and B(103)) xor (A(56) and B(102)) xor (A(57) and B(101)) xor (A(58) and B(100)) xor (A(59) and B(99)) xor (A(60) and B(98)) xor (A(61) and B(97)) xor (A(62) and B(96)) xor (A(63) and B(95)) xor (A(64) and B(94)) xor (A(65) and B(93)) xor (A(66) and B(92)) xor (A(67) and B(91)) xor (A(68) and B(90)) xor (A(69) and B(89)) xor (A(70) and B(88)) xor (A(71) and B(87)) xor (A(72) and B(86)) xor (A(73) and B(85)) xor (A(74) and B(84)) xor (A(75) and B(83)) xor (A(76) and B(82)) xor (A(77) and B(81)) xor (A(78) and B(80)) xor (A(79) and B(79)) xor (A(80) and B(78)) xor (A(81) and B(77)) xor (A(82) and B(76)) xor (A(83) and B(75)) xor (A(84) and B(74)) xor (A(85) and B(73)) xor (A(86) and B(72)) xor (A(87) and B(71)) xor (A(88) and B(70)) xor (A(89) and B(69)) xor (A(90) and B(68)) xor (A(91) and B(67)) xor (A(92) and B(66)) xor (A(93) and B(65)) xor (A(94) and B(64)) xor (A(95) and B(63)) xor (A(96) and B(62)) xor (A(97) and B(61)) xor (A(98) and B(60)) xor (A(99) and B(59)) xor (A(100) and B(58)) xor (A(101) and B(57)) xor (A(102) and B(56)) xor (A(103) and B(55)) xor (A(104) and B(54)) xor (A(105) and B(53)) xor (A(106) and B(52)) xor (A(107) and B(51)) xor (A(108) and B(50)) xor (A(109) and B(49)) xor (A(110) and B(48)) xor (A(111) and B(47)) xor (A(112) and B(46)) xor (A(113) and B(45)) xor (A(114) and B(44)) xor (A(115) and B(43)) xor (A(116) and B(42)) xor (A(117) and B(41)) xor (A(118) and B(40)) xor (A(119) and B(39)) xor (A(120) and B(38)) xor (A(121) and B(37)) xor (A(122) and B(36)) xor (A(123) and B(35)) xor (A(124) and B(34)) xor (A(125) and B(33)) xor (A(126) and B(32)) xor (A(36) and B(127)) xor (A(37) and B(126)) xor (A(38) and B(125)) xor (A(39) and B(124)) xor (A(40) and B(123)) xor (A(41) and B(122)) xor (A(42) and B(121)) xor (A(43) and B(120)) xor (A(44) and B(119)) xor (A(45) and B(118)) xor (A(46) and B(117)) xor (A(47) and B(116)) xor (A(48) and B(115)) xor (A(49) and B(114)) xor (A(50) and B(113)) xor (A(51) and B(112)) xor (A(52) and B(111)) xor (A(53) and B(110)) xor (A(54) and B(109)) xor (A(55) and B(108)) xor (A(56) and B(107)) xor (A(57) and B(106)) xor (A(58) and B(105)) xor (A(59) and B(104)) xor (A(60) and B(103)) xor (A(61) and B(102)) xor (A(62) and B(101)) xor (A(63) and B(100)) xor (A(64) and B(99)) xor (A(65) and B(98)) xor (A(66) and B(97)) xor (A(67) and B(96)) xor (A(68) and B(95)) xor (A(69) and B(94)) xor (A(70) and B(93)) xor (A(71) and B(92)) xor (A(72) and B(91)) xor (A(73) and B(90)) xor (A(74) and B(89)) xor (A(75) and B(88)) xor (A(76) and B(87)) xor (A(77) and B(86)) xor (A(78) and B(85)) xor (A(79) and B(84)) xor (A(80) and B(83)) xor (A(81) and B(82)) xor (A(82) and B(81)) xor (A(83) and B(80)) xor (A(84) and B(79)) xor (A(85) and B(78)) xor (A(86) and B(77)) xor (A(87) and B(76)) xor (A(88) and B(75)) xor (A(89) and B(74)) xor (A(90) and B(73)) xor (A(91) and B(72)) xor (A(92) and B(71)) xor (A(93) and B(70)) xor (A(94) and B(69)) xor (A(95) and B(68)) xor (A(96) and B(67)) xor (A(97) and B(66)) xor (A(98) and B(65)) xor (A(99) and B(64)) xor (A(100) and B(63)) xor (A(101) and B(62)) xor (A(102) and B(61)) xor (A(103) and B(60)) xor (A(104) and B(59)) xor (A(105) and B(58)) xor (A(106) and B(57)) xor (A(107) and B(56)) xor (A(108) and B(55)) xor (A(109) and B(54)) xor (A(110) and B(53)) xor (A(111) and B(52)) xor (A(112) and B(51)) xor (A(113) and B(50)) xor (A(114) and B(49)) xor (A(115) and B(48)) xor (A(116) and B(47)) xor (A(117) and B(46)) xor (A(118) and B(45)) xor (A(119) and B(44)) xor (A(120) and B(43)) xor (A(121) and B(42)) xor (A(122) and B(41)) xor (A(123) and B(40)) xor (A(124) and B(39)) xor (A(125) and B(38)) xor (A(126) and B(37)) xor (A(37) and B(127)) xor (A(38) and B(126)) xor (A(39) and B(125)) xor (A(40) and B(124)) xor (A(41) and B(123)) xor (A(42) and B(122)) xor (A(43) and B(121)) xor (A(44) and B(120)) xor (A(45) and B(119)) xor (A(46) and B(118)) xor (A(47) and B(117)) xor (A(48) and B(116)) xor (A(49) and B(115)) xor (A(50) and B(114)) xor (A(51) and B(113)) xor (A(52) and B(112)) xor (A(53) and B(111)) xor (A(54) and B(110)) xor (A(55) and B(109)) xor (A(56) and B(108)) xor (A(57) and B(107)) xor (A(58) and B(106)) xor (A(59) and B(105)) xor (A(60) and B(104)) xor (A(61) and B(103)) xor (A(62) and B(102)) xor (A(63) and B(101)) xor (A(64) and B(100)) xor (A(65) and B(99)) xor (A(66) and B(98)) xor (A(67) and B(97)) xor (A(68) and B(96)) xor (A(69) and B(95)) xor (A(70) and B(94)) xor (A(71) and B(93)) xor (A(72) and B(92)) xor (A(73) and B(91)) xor (A(74) and B(90)) xor (A(75) and B(89)) xor (A(76) and B(88)) xor (A(77) and B(87)) xor (A(78) and B(86)) xor (A(79) and B(85)) xor (A(80) and B(84)) xor (A(81) and B(83)) xor (A(82) and B(82)) xor (A(83) and B(81)) xor (A(84) and B(80)) xor (A(85) and B(79)) xor (A(86) and B(78)) xor (A(87) and B(77)) xor (A(88) and B(76)) xor (A(89) and B(75)) xor (A(90) and B(74)) xor (A(91) and B(73)) xor (A(92) and B(72)) xor (A(93) and B(71)) xor (A(94) and B(70)) xor (A(95) and B(69)) xor (A(96) and B(68)) xor (A(97) and B(67)) xor (A(98) and B(66)) xor (A(99) and B(65)) xor (A(100) and B(64)) xor (A(101) and B(63)) xor (A(102) and B(62)) xor (A(103) and B(61)) xor (A(104) and B(60)) xor (A(105) and B(59)) xor (A(106) and B(58)) xor (A(107) and B(57)) xor (A(108) and B(56)) xor (A(109) and B(55)) xor (A(110) and B(54)) xor (A(111) and B(53)) xor (A(112) and B(52)) xor (A(113) and B(51)) xor (A(114) and B(50)) xor (A(115) and B(49)) xor (A(116) and B(48)) xor (A(117) and B(47)) xor (A(118) and B(46)) xor (A(119) and B(45)) xor (A(120) and B(44)) xor (A(121) and B(43)) xor (A(122) and B(42)) xor (A(123) and B(41)) xor (A(124) and B(40)) xor (A(125) and B(39)) xor (A(126) and B(38)) xor (A(38) and B(127)) xor (A(39) and B(126)) xor (A(40) and B(125)) xor (A(41) and B(124)) xor (A(42) and B(123)) xor (A(43) and B(122)) xor (A(44) and B(121)) xor (A(45) and B(120)) xor (A(46) and B(119)) xor (A(47) and B(118)) xor (A(48) and B(117)) xor (A(49) and B(116)) xor (A(50) and B(115)) xor (A(51) and B(114)) xor (A(52) and B(113)) xor (A(53) and B(112)) xor (A(54) and B(111)) xor (A(55) and B(110)) xor (A(56) and B(109)) xor (A(57) and B(108)) xor (A(58) and B(107)) xor (A(59) and B(106)) xor (A(60) and B(105)) xor (A(61) and B(104)) xor (A(62) and B(103)) xor (A(63) and B(102)) xor (A(64) and B(101)) xor (A(65) and B(100)) xor (A(66) and B(99)) xor (A(67) and B(98)) xor (A(68) and B(97)) xor (A(69) and B(96)) xor (A(70) and B(95)) xor (A(71) and B(94)) xor (A(72) and B(93)) xor (A(73) and B(92)) xor (A(74) and B(91)) xor (A(75) and B(90)) xor (A(76) and B(89)) xor (A(77) and B(88)) xor (A(78) and B(87)) xor (A(79) and B(86)) xor (A(80) and B(85)) xor (A(81) and B(84)) xor (A(82) and B(83)) xor (A(83) and B(82)) xor (A(84) and B(81)) xor (A(85) and B(80)) xor (A(86) and B(79)) xor (A(87) and B(78)) xor (A(88) and B(77)) xor (A(89) and B(76)) xor (A(90) and B(75)) xor (A(91) and B(74)) xor (A(92) and B(73)) xor (A(93) and B(72)) xor (A(94) and B(71)) xor (A(95) and B(70)) xor (A(96) and B(69)) xor (A(97) and B(68)) xor (A(98) and B(67)) xor (A(99) and B(66)) xor (A(100) and B(65)) xor (A(101) and B(64)) xor (A(102) and B(63)) xor (A(103) and B(62)) xor (A(104) and B(61)) xor (A(105) and B(60)) xor (A(106) and B(59)) xor (A(107) and B(58)) xor (A(108) and B(57)) xor (A(109) and B(56)) xor (A(110) and B(55)) xor (A(111) and B(54)) xor (A(112) and B(53)) xor (A(113) and B(52)) xor (A(114) and B(51)) xor (A(115) and B(50)) xor (A(116) and B(49)) xor (A(117) and B(48)) xor (A(118) and B(47)) xor (A(119) and B(46)) xor (A(120) and B(45)) xor (A(121) and B(44)) xor (A(122) and B(43)) xor (A(123) and B(42)) xor (A(124) and B(41)) xor (A(125) and B(40)) xor (A(126) and B(40));
    C(39)  <= (A(0) and B(39)) xor (A(1) and B(38)) xor (A(2) and B(37)) xor (A(3) and B(36)) xor (A(4) and B(35)) xor (A(5) and B(34)) xor (A(6) and B(33)) xor (A(7) and B(32)) xor (A(8) and B(31)) xor (A(9) and B(30)) xor (A(10) and B(29)) xor (A(11) and B(28)) xor (A(12) and B(27)) xor (A(13) and B(26)) xor (A(14) and B(25)) xor (A(15) and B(24)) xor (A(16) and B(23)) xor (A(17) and B(23)) xor (A(18) and B(21)) xor (A(19) and B(20)) xor (A(20) and B(19)) xor (A(21) and B(18)) xor (A(23) and B(17)) xor (A(23) and B(16)) xor (A(24) and B(15)) xor (A(25) and B(14)) xor (A(26) and B(13)) xor (A(27) and B(12)) xor (A(28) and B(11)) xor (A(29) and B(10)) xor (A(30) and B(9)) xor (A(31) and B(8)) xor (A(32) and B(7)) xor (A(33) and B(6)) xor (A(34) and B(5)) xor (A(35) and B(4)) xor (A(36) and B(3)) xor (A(37) and B(2)) xor (A(38) and B(1)) xor (A(39) and B(0)) xor (A(32) and B(127)) xor (A(33) and B(126)) xor (A(34) and B(125)) xor (A(35) and B(124)) xor (A(36) and B(123)) xor (A(37) and B(122)) xor (A(38) and B(121)) xor (A(39) and B(120)) xor (A(40) and B(119)) xor (A(41) and B(118)) xor (A(42) and B(117)) xor (A(43) and B(116)) xor (A(44) and B(115)) xor (A(45) and B(114)) xor (A(46) and B(113)) xor (A(47) and B(112)) xor (A(48) and B(111)) xor (A(49) and B(110)) xor (A(50) and B(109)) xor (A(51) and B(108)) xor (A(52) and B(107)) xor (A(53) and B(106)) xor (A(54) and B(105)) xor (A(55) and B(104)) xor (A(56) and B(103)) xor (A(57) and B(102)) xor (A(58) and B(101)) xor (A(59) and B(100)) xor (A(60) and B(99)) xor (A(61) and B(98)) xor (A(62) and B(97)) xor (A(63) and B(96)) xor (A(64) and B(95)) xor (A(65) and B(94)) xor (A(66) and B(93)) xor (A(67) and B(92)) xor (A(68) and B(91)) xor (A(69) and B(90)) xor (A(70) and B(89)) xor (A(71) and B(88)) xor (A(72) and B(87)) xor (A(73) and B(86)) xor (A(74) and B(85)) xor (A(75) and B(84)) xor (A(76) and B(83)) xor (A(77) and B(82)) xor (A(78) and B(81)) xor (A(79) and B(80)) xor (A(80) and B(79)) xor (A(81) and B(78)) xor (A(82) and B(77)) xor (A(83) and B(76)) xor (A(84) and B(75)) xor (A(85) and B(74)) xor (A(86) and B(73)) xor (A(87) and B(72)) xor (A(88) and B(71)) xor (A(89) and B(70)) xor (A(90) and B(69)) xor (A(91) and B(68)) xor (A(92) and B(67)) xor (A(93) and B(66)) xor (A(94) and B(65)) xor (A(95) and B(64)) xor (A(96) and B(63)) xor (A(97) and B(62)) xor (A(98) and B(61)) xor (A(99) and B(60)) xor (A(100) and B(59)) xor (A(101) and B(58)) xor (A(102) and B(57)) xor (A(103) and B(56)) xor (A(104) and B(55)) xor (A(105) and B(54)) xor (A(106) and B(53)) xor (A(107) and B(52)) xor (A(108) and B(51)) xor (A(109) and B(50)) xor (A(110) and B(49)) xor (A(111) and B(48)) xor (A(112) and B(47)) xor (A(113) and B(46)) xor (A(114) and B(45)) xor (A(115) and B(44)) xor (A(116) and B(43)) xor (A(117) and B(42)) xor (A(118) and B(41)) xor (A(119) and B(40)) xor (A(120) and B(39)) xor (A(121) and B(38)) xor (A(122) and B(37)) xor (A(123) and B(36)) xor (A(124) and B(35)) xor (A(125) and B(34)) xor (A(126) and B(33)) xor (A(37) and B(127)) xor (A(38) and B(126)) xor (A(39) and B(125)) xor (A(40) and B(124)) xor (A(41) and B(123)) xor (A(42) and B(122)) xor (A(43) and B(121)) xor (A(44) and B(120)) xor (A(45) and B(119)) xor (A(46) and B(118)) xor (A(47) and B(117)) xor (A(48) and B(116)) xor (A(49) and B(115)) xor (A(50) and B(114)) xor (A(51) and B(113)) xor (A(52) and B(112)) xor (A(53) and B(111)) xor (A(54) and B(110)) xor (A(55) and B(109)) xor (A(56) and B(108)) xor (A(57) and B(107)) xor (A(58) and B(106)) xor (A(59) and B(105)) xor (A(60) and B(104)) xor (A(61) and B(103)) xor (A(62) and B(102)) xor (A(63) and B(101)) xor (A(64) and B(100)) xor (A(65) and B(99)) xor (A(66) and B(98)) xor (A(67) and B(97)) xor (A(68) and B(96)) xor (A(69) and B(95)) xor (A(70) and B(94)) xor (A(71) and B(93)) xor (A(72) and B(92)) xor (A(73) and B(91)) xor (A(74) and B(90)) xor (A(75) and B(89)) xor (A(76) and B(88)) xor (A(77) and B(87)) xor (A(78) and B(86)) xor (A(79) and B(85)) xor (A(80) and B(84)) xor (A(81) and B(83)) xor (A(82) and B(82)) xor (A(83) and B(81)) xor (A(84) and B(80)) xor (A(85) and B(79)) xor (A(86) and B(78)) xor (A(87) and B(77)) xor (A(88) and B(76)) xor (A(89) and B(75)) xor (A(90) and B(74)) xor (A(91) and B(73)) xor (A(92) and B(72)) xor (A(93) and B(71)) xor (A(94) and B(70)) xor (A(95) and B(69)) xor (A(96) and B(68)) xor (A(97) and B(67)) xor (A(98) and B(66)) xor (A(99) and B(65)) xor (A(100) and B(64)) xor (A(101) and B(63)) xor (A(102) and B(62)) xor (A(103) and B(61)) xor (A(104) and B(60)) xor (A(105) and B(59)) xor (A(106) and B(58)) xor (A(107) and B(57)) xor (A(108) and B(56)) xor (A(109) and B(55)) xor (A(110) and B(54)) xor (A(111) and B(53)) xor (A(112) and B(52)) xor (A(113) and B(51)) xor (A(114) and B(50)) xor (A(115) and B(49)) xor (A(116) and B(48)) xor (A(117) and B(47)) xor (A(118) and B(46)) xor (A(119) and B(45)) xor (A(120) and B(44)) xor (A(121) and B(43)) xor (A(122) and B(42)) xor (A(123) and B(41)) xor (A(124) and B(40)) xor (A(125) and B(39)) xor (A(126) and B(38)) xor (A(38) and B(127)) xor (A(39) and B(126)) xor (A(40) and B(125)) xor (A(41) and B(124)) xor (A(42) and B(123)) xor (A(43) and B(122)) xor (A(44) and B(121)) xor (A(45) and B(120)) xor (A(46) and B(119)) xor (A(47) and B(118)) xor (A(48) and B(117)) xor (A(49) and B(116)) xor (A(50) and B(115)) xor (A(51) and B(114)) xor (A(52) and B(113)) xor (A(53) and B(112)) xor (A(54) and B(111)) xor (A(55) and B(110)) xor (A(56) and B(109)) xor (A(57) and B(108)) xor (A(58) and B(107)) xor (A(59) and B(106)) xor (A(60) and B(105)) xor (A(61) and B(104)) xor (A(62) and B(103)) xor (A(63) and B(102)) xor (A(64) and B(101)) xor (A(65) and B(100)) xor (A(66) and B(99)) xor (A(67) and B(98)) xor (A(68) and B(97)) xor (A(69) and B(96)) xor (A(70) and B(95)) xor (A(71) and B(94)) xor (A(72) and B(93)) xor (A(73) and B(92)) xor (A(74) and B(91)) xor (A(75) and B(90)) xor (A(76) and B(89)) xor (A(77) and B(88)) xor (A(78) and B(87)) xor (A(79) and B(86)) xor (A(80) and B(85)) xor (A(81) and B(84)) xor (A(82) and B(83)) xor (A(83) and B(82)) xor (A(84) and B(81)) xor (A(85) and B(80)) xor (A(86) and B(79)) xor (A(87) and B(78)) xor (A(88) and B(77)) xor (A(89) and B(76)) xor (A(90) and B(75)) xor (A(91) and B(74)) xor (A(92) and B(73)) xor (A(93) and B(72)) xor (A(94) and B(71)) xor (A(95) and B(70)) xor (A(96) and B(69)) xor (A(97) and B(68)) xor (A(98) and B(67)) xor (A(99) and B(66)) xor (A(100) and B(65)) xor (A(101) and B(64)) xor (A(102) and B(63)) xor (A(103) and B(62)) xor (A(104) and B(61)) xor (A(105) and B(60)) xor (A(106) and B(59)) xor (A(107) and B(58)) xor (A(108) and B(57)) xor (A(109) and B(56)) xor (A(110) and B(55)) xor (A(111) and B(54)) xor (A(112) and B(53)) xor (A(113) and B(52)) xor (A(114) and B(51)) xor (A(115) and B(50)) xor (A(116) and B(49)) xor (A(117) and B(48)) xor (A(118) and B(47)) xor (A(119) and B(46)) xor (A(120) and B(45)) xor (A(121) and B(44)) xor (A(122) and B(43)) xor (A(123) and B(42)) xor (A(124) and B(41)) xor (A(125) and B(40)) xor (A(126) and B(39)) xor (A(39) and B(127)) xor (A(40) and B(126)) xor (A(41) and B(125)) xor (A(42) and B(124)) xor (A(43) and B(123)) xor (A(44) and B(122)) xor (A(45) and B(121)) xor (A(46) and B(120)) xor (A(47) and B(119)) xor (A(48) and B(118)) xor (A(49) and B(117)) xor (A(50) and B(116)) xor (A(51) and B(115)) xor (A(52) and B(114)) xor (A(53) and B(113)) xor (A(54) and B(112)) xor (A(55) and B(111)) xor (A(56) and B(110)) xor (A(57) and B(109)) xor (A(58) and B(108)) xor (A(59) and B(107)) xor (A(60) and B(106)) xor (A(61) and B(105)) xor (A(62) and B(104)) xor (A(63) and B(103)) xor (A(64) and B(102)) xor (A(65) and B(101)) xor (A(66) and B(100)) xor (A(67) and B(99)) xor (A(68) and B(98)) xor (A(69) and B(97)) xor (A(70) and B(96)) xor (A(71) and B(95)) xor (A(72) and B(94)) xor (A(73) and B(93)) xor (A(74) and B(92)) xor (A(75) and B(91)) xor (A(76) and B(90)) xor (A(77) and B(89)) xor (A(78) and B(88)) xor (A(79) and B(87)) xor (A(80) and B(86)) xor (A(81) and B(85)) xor (A(82) and B(84)) xor (A(83) and B(83)) xor (A(84) and B(82)) xor (A(85) and B(81)) xor (A(86) and B(80)) xor (A(87) and B(79)) xor (A(88) and B(78)) xor (A(89) and B(77)) xor (A(90) and B(76)) xor (A(91) and B(75)) xor (A(92) and B(74)) xor (A(93) and B(73)) xor (A(94) and B(72)) xor (A(95) and B(71)) xor (A(96) and B(70)) xor (A(97) and B(69)) xor (A(98) and B(68)) xor (A(99) and B(67)) xor (A(100) and B(66)) xor (A(101) and B(65)) xor (A(102) and B(64)) xor (A(103) and B(63)) xor (A(104) and B(62)) xor (A(105) and B(61)) xor (A(106) and B(60)) xor (A(107) and B(59)) xor (A(108) and B(58)) xor (A(109) and B(57)) xor (A(110) and B(56)) xor (A(111) and B(55)) xor (A(112) and B(54)) xor (A(113) and B(53)) xor (A(114) and B(52)) xor (A(115) and B(51)) xor (A(116) and B(50)) xor (A(117) and B(49)) xor (A(118) and B(48)) xor (A(119) and B(47)) xor (A(120) and B(46)) xor (A(121) and B(45)) xor (A(122) and B(44)) xor (A(123) and B(43)) xor (A(124) and B(42)) xor (A(125) and B(41)) xor (A(126) and B(41));
    C(40)  <= (A(0) and B(40)) xor (A(1) and B(39)) xor (A(2) and B(38)) xor (A(3) and B(37)) xor (A(4) and B(36)) xor (A(5) and B(35)) xor (A(6) and B(34)) xor (A(7) and B(33)) xor (A(8) and B(32)) xor (A(9) and B(31)) xor (A(10) and B(30)) xor (A(11) and B(29)) xor (A(12) and B(28)) xor (A(13) and B(27)) xor (A(14) and B(26)) xor (A(15) and B(25)) xor (A(16) and B(24)) xor (A(17) and B(23)) xor (A(18) and B(23)) xor (A(19) and B(21)) xor (A(20) and B(20)) xor (A(21) and B(19)) xor (A(23) and B(18)) xor (A(23) and B(17)) xor (A(24) and B(16)) xor (A(25) and B(15)) xor (A(26) and B(14)) xor (A(27) and B(13)) xor (A(28) and B(12)) xor (A(29) and B(11)) xor (A(30) and B(10)) xor (A(31) and B(9)) xor (A(32) and B(8)) xor (A(33) and B(7)) xor (A(34) and B(6)) xor (A(35) and B(5)) xor (A(36) and B(4)) xor (A(37) and B(3)) xor (A(38) and B(2)) xor (A(39) and B(1)) xor (A(40) and B(0)) xor (A(33) and B(127)) xor (A(34) and B(126)) xor (A(35) and B(125)) xor (A(36) and B(124)) xor (A(37) and B(123)) xor (A(38) and B(122)) xor (A(39) and B(121)) xor (A(40) and B(120)) xor (A(41) and B(119)) xor (A(42) and B(118)) xor (A(43) and B(117)) xor (A(44) and B(116)) xor (A(45) and B(115)) xor (A(46) and B(114)) xor (A(47) and B(113)) xor (A(48) and B(112)) xor (A(49) and B(111)) xor (A(50) and B(110)) xor (A(51) and B(109)) xor (A(52) and B(108)) xor (A(53) and B(107)) xor (A(54) and B(106)) xor (A(55) and B(105)) xor (A(56) and B(104)) xor (A(57) and B(103)) xor (A(58) and B(102)) xor (A(59) and B(101)) xor (A(60) and B(100)) xor (A(61) and B(99)) xor (A(62) and B(98)) xor (A(63) and B(97)) xor (A(64) and B(96)) xor (A(65) and B(95)) xor (A(66) and B(94)) xor (A(67) and B(93)) xor (A(68) and B(92)) xor (A(69) and B(91)) xor (A(70) and B(90)) xor (A(71) and B(89)) xor (A(72) and B(88)) xor (A(73) and B(87)) xor (A(74) and B(86)) xor (A(75) and B(85)) xor (A(76) and B(84)) xor (A(77) and B(83)) xor (A(78) and B(82)) xor (A(79) and B(81)) xor (A(80) and B(80)) xor (A(81) and B(79)) xor (A(82) and B(78)) xor (A(83) and B(77)) xor (A(84) and B(76)) xor (A(85) and B(75)) xor (A(86) and B(74)) xor (A(87) and B(73)) xor (A(88) and B(72)) xor (A(89) and B(71)) xor (A(90) and B(70)) xor (A(91) and B(69)) xor (A(92) and B(68)) xor (A(93) and B(67)) xor (A(94) and B(66)) xor (A(95) and B(65)) xor (A(96) and B(64)) xor (A(97) and B(63)) xor (A(98) and B(62)) xor (A(99) and B(61)) xor (A(100) and B(60)) xor (A(101) and B(59)) xor (A(102) and B(58)) xor (A(103) and B(57)) xor (A(104) and B(56)) xor (A(105) and B(55)) xor (A(106) and B(54)) xor (A(107) and B(53)) xor (A(108) and B(52)) xor (A(109) and B(51)) xor (A(110) and B(50)) xor (A(111) and B(49)) xor (A(112) and B(48)) xor (A(113) and B(47)) xor (A(114) and B(46)) xor (A(115) and B(45)) xor (A(116) and B(44)) xor (A(117) and B(43)) xor (A(118) and B(42)) xor (A(119) and B(41)) xor (A(120) and B(40)) xor (A(121) and B(39)) xor (A(122) and B(38)) xor (A(123) and B(37)) xor (A(124) and B(36)) xor (A(125) and B(35)) xor (A(126) and B(34)) xor (A(38) and B(127)) xor (A(39) and B(126)) xor (A(40) and B(125)) xor (A(41) and B(124)) xor (A(42) and B(123)) xor (A(43) and B(122)) xor (A(44) and B(121)) xor (A(45) and B(120)) xor (A(46) and B(119)) xor (A(47) and B(118)) xor (A(48) and B(117)) xor (A(49) and B(116)) xor (A(50) and B(115)) xor (A(51) and B(114)) xor (A(52) and B(113)) xor (A(53) and B(112)) xor (A(54) and B(111)) xor (A(55) and B(110)) xor (A(56) and B(109)) xor (A(57) and B(108)) xor (A(58) and B(107)) xor (A(59) and B(106)) xor (A(60) and B(105)) xor (A(61) and B(104)) xor (A(62) and B(103)) xor (A(63) and B(102)) xor (A(64) and B(101)) xor (A(65) and B(100)) xor (A(66) and B(99)) xor (A(67) and B(98)) xor (A(68) and B(97)) xor (A(69) and B(96)) xor (A(70) and B(95)) xor (A(71) and B(94)) xor (A(72) and B(93)) xor (A(73) and B(92)) xor (A(74) and B(91)) xor (A(75) and B(90)) xor (A(76) and B(89)) xor (A(77) and B(88)) xor (A(78) and B(87)) xor (A(79) and B(86)) xor (A(80) and B(85)) xor (A(81) and B(84)) xor (A(82) and B(83)) xor (A(83) and B(82)) xor (A(84) and B(81)) xor (A(85) and B(80)) xor (A(86) and B(79)) xor (A(87) and B(78)) xor (A(88) and B(77)) xor (A(89) and B(76)) xor (A(90) and B(75)) xor (A(91) and B(74)) xor (A(92) and B(73)) xor (A(93) and B(72)) xor (A(94) and B(71)) xor (A(95) and B(70)) xor (A(96) and B(69)) xor (A(97) and B(68)) xor (A(98) and B(67)) xor (A(99) and B(66)) xor (A(100) and B(65)) xor (A(101) and B(64)) xor (A(102) and B(63)) xor (A(103) and B(62)) xor (A(104) and B(61)) xor (A(105) and B(60)) xor (A(106) and B(59)) xor (A(107) and B(58)) xor (A(108) and B(57)) xor (A(109) and B(56)) xor (A(110) and B(55)) xor (A(111) and B(54)) xor (A(112) and B(53)) xor (A(113) and B(52)) xor (A(114) and B(51)) xor (A(115) and B(50)) xor (A(116) and B(49)) xor (A(117) and B(48)) xor (A(118) and B(47)) xor (A(119) and B(46)) xor (A(120) and B(45)) xor (A(121) and B(44)) xor (A(122) and B(43)) xor (A(123) and B(42)) xor (A(124) and B(41)) xor (A(125) and B(40)) xor (A(126) and B(39)) xor (A(39) and B(127)) xor (A(40) and B(126)) xor (A(41) and B(125)) xor (A(42) and B(124)) xor (A(43) and B(123)) xor (A(44) and B(122)) xor (A(45) and B(121)) xor (A(46) and B(120)) xor (A(47) and B(119)) xor (A(48) and B(118)) xor (A(49) and B(117)) xor (A(50) and B(116)) xor (A(51) and B(115)) xor (A(52) and B(114)) xor (A(53) and B(113)) xor (A(54) and B(112)) xor (A(55) and B(111)) xor (A(56) and B(110)) xor (A(57) and B(109)) xor (A(58) and B(108)) xor (A(59) and B(107)) xor (A(60) and B(106)) xor (A(61) and B(105)) xor (A(62) and B(104)) xor (A(63) and B(103)) xor (A(64) and B(102)) xor (A(65) and B(101)) xor (A(66) and B(100)) xor (A(67) and B(99)) xor (A(68) and B(98)) xor (A(69) and B(97)) xor (A(70) and B(96)) xor (A(71) and B(95)) xor (A(72) and B(94)) xor (A(73) and B(93)) xor (A(74) and B(92)) xor (A(75) and B(91)) xor (A(76) and B(90)) xor (A(77) and B(89)) xor (A(78) and B(88)) xor (A(79) and B(87)) xor (A(80) and B(86)) xor (A(81) and B(85)) xor (A(82) and B(84)) xor (A(83) and B(83)) xor (A(84) and B(82)) xor (A(85) and B(81)) xor (A(86) and B(80)) xor (A(87) and B(79)) xor (A(88) and B(78)) xor (A(89) and B(77)) xor (A(90) and B(76)) xor (A(91) and B(75)) xor (A(92) and B(74)) xor (A(93) and B(73)) xor (A(94) and B(72)) xor (A(95) and B(71)) xor (A(96) and B(70)) xor (A(97) and B(69)) xor (A(98) and B(68)) xor (A(99) and B(67)) xor (A(100) and B(66)) xor (A(101) and B(65)) xor (A(102) and B(64)) xor (A(103) and B(63)) xor (A(104) and B(62)) xor (A(105) and B(61)) xor (A(106) and B(60)) xor (A(107) and B(59)) xor (A(108) and B(58)) xor (A(109) and B(57)) xor (A(110) and B(56)) xor (A(111) and B(55)) xor (A(112) and B(54)) xor (A(113) and B(53)) xor (A(114) and B(52)) xor (A(115) and B(51)) xor (A(116) and B(50)) xor (A(117) and B(49)) xor (A(118) and B(48)) xor (A(119) and B(47)) xor (A(120) and B(46)) xor (A(121) and B(45)) xor (A(122) and B(44)) xor (A(123) and B(43)) xor (A(124) and B(42)) xor (A(125) and B(41)) xor (A(126) and B(40)) xor (A(40) and B(127)) xor (A(41) and B(126)) xor (A(42) and B(125)) xor (A(43) and B(124)) xor (A(44) and B(123)) xor (A(45) and B(122)) xor (A(46) and B(121)) xor (A(47) and B(120)) xor (A(48) and B(119)) xor (A(49) and B(118)) xor (A(50) and B(117)) xor (A(51) and B(116)) xor (A(52) and B(115)) xor (A(53) and B(114)) xor (A(54) and B(113)) xor (A(55) and B(112)) xor (A(56) and B(111)) xor (A(57) and B(110)) xor (A(58) and B(109)) xor (A(59) and B(108)) xor (A(60) and B(107)) xor (A(61) and B(106)) xor (A(62) and B(105)) xor (A(63) and B(104)) xor (A(64) and B(103)) xor (A(65) and B(102)) xor (A(66) and B(101)) xor (A(67) and B(100)) xor (A(68) and B(99)) xor (A(69) and B(98)) xor (A(70) and B(97)) xor (A(71) and B(96)) xor (A(72) and B(95)) xor (A(73) and B(94)) xor (A(74) and B(93)) xor (A(75) and B(92)) xor (A(76) and B(91)) xor (A(77) and B(90)) xor (A(78) and B(89)) xor (A(79) and B(88)) xor (A(80) and B(87)) xor (A(81) and B(86)) xor (A(82) and B(85)) xor (A(83) and B(84)) xor (A(84) and B(83)) xor (A(85) and B(82)) xor (A(86) and B(81)) xor (A(87) and B(80)) xor (A(88) and B(79)) xor (A(89) and B(78)) xor (A(90) and B(77)) xor (A(91) and B(76)) xor (A(92) and B(75)) xor (A(93) and B(74)) xor (A(94) and B(73)) xor (A(95) and B(72)) xor (A(96) and B(71)) xor (A(97) and B(70)) xor (A(98) and B(69)) xor (A(99) and B(68)) xor (A(100) and B(67)) xor (A(101) and B(66)) xor (A(102) and B(65)) xor (A(103) and B(64)) xor (A(104) and B(63)) xor (A(105) and B(62)) xor (A(106) and B(61)) xor (A(107) and B(60)) xor (A(108) and B(59)) xor (A(109) and B(58)) xor (A(110) and B(57)) xor (A(111) and B(56)) xor (A(112) and B(55)) xor (A(113) and B(54)) xor (A(114) and B(53)) xor (A(115) and B(52)) xor (A(116) and B(51)) xor (A(117) and B(50)) xor (A(118) and B(49)) xor (A(119) and B(48)) xor (A(120) and B(47)) xor (A(121) and B(46)) xor (A(122) and B(45)) xor (A(123) and B(44)) xor (A(124) and B(43)) xor (A(125) and B(42)) xor (A(126) and B(42));
    C(41)  <= (A(0) and B(41)) xor (A(1) and B(40)) xor (A(2) and B(39)) xor (A(3) and B(38)) xor (A(4) and B(37)) xor (A(5) and B(36)) xor (A(6) and B(35)) xor (A(7) and B(34)) xor (A(8) and B(33)) xor (A(9) and B(32)) xor (A(10) and B(31)) xor (A(11) and B(30)) xor (A(12) and B(29)) xor (A(13) and B(28)) xor (A(14) and B(27)) xor (A(15) and B(26)) xor (A(16) and B(25)) xor (A(17) and B(24)) xor (A(18) and B(23)) xor (A(19) and B(23)) xor (A(20) and B(21)) xor (A(21) and B(20)) xor (A(23) and B(19)) xor (A(23) and B(18)) xor (A(24) and B(17)) xor (A(25) and B(16)) xor (A(26) and B(15)) xor (A(27) and B(14)) xor (A(28) and B(13)) xor (A(29) and B(12)) xor (A(30) and B(11)) xor (A(31) and B(10)) xor (A(32) and B(9)) xor (A(33) and B(8)) xor (A(34) and B(7)) xor (A(35) and B(6)) xor (A(36) and B(5)) xor (A(37) and B(4)) xor (A(38) and B(3)) xor (A(39) and B(2)) xor (A(40) and B(1)) xor (A(41) and B(0)) xor (A(34) and B(127)) xor (A(35) and B(126)) xor (A(36) and B(125)) xor (A(37) and B(124)) xor (A(38) and B(123)) xor (A(39) and B(122)) xor (A(40) and B(121)) xor (A(41) and B(120)) xor (A(42) and B(119)) xor (A(43) and B(118)) xor (A(44) and B(117)) xor (A(45) and B(116)) xor (A(46) and B(115)) xor (A(47) and B(114)) xor (A(48) and B(113)) xor (A(49) and B(112)) xor (A(50) and B(111)) xor (A(51) and B(110)) xor (A(52) and B(109)) xor (A(53) and B(108)) xor (A(54) and B(107)) xor (A(55) and B(106)) xor (A(56) and B(105)) xor (A(57) and B(104)) xor (A(58) and B(103)) xor (A(59) and B(102)) xor (A(60) and B(101)) xor (A(61) and B(100)) xor (A(62) and B(99)) xor (A(63) and B(98)) xor (A(64) and B(97)) xor (A(65) and B(96)) xor (A(66) and B(95)) xor (A(67) and B(94)) xor (A(68) and B(93)) xor (A(69) and B(92)) xor (A(70) and B(91)) xor (A(71) and B(90)) xor (A(72) and B(89)) xor (A(73) and B(88)) xor (A(74) and B(87)) xor (A(75) and B(86)) xor (A(76) and B(85)) xor (A(77) and B(84)) xor (A(78) and B(83)) xor (A(79) and B(82)) xor (A(80) and B(81)) xor (A(81) and B(80)) xor (A(82) and B(79)) xor (A(83) and B(78)) xor (A(84) and B(77)) xor (A(85) and B(76)) xor (A(86) and B(75)) xor (A(87) and B(74)) xor (A(88) and B(73)) xor (A(89) and B(72)) xor (A(90) and B(71)) xor (A(91) and B(70)) xor (A(92) and B(69)) xor (A(93) and B(68)) xor (A(94) and B(67)) xor (A(95) and B(66)) xor (A(96) and B(65)) xor (A(97) and B(64)) xor (A(98) and B(63)) xor (A(99) and B(62)) xor (A(100) and B(61)) xor (A(101) and B(60)) xor (A(102) and B(59)) xor (A(103) and B(58)) xor (A(104) and B(57)) xor (A(105) and B(56)) xor (A(106) and B(55)) xor (A(107) and B(54)) xor (A(108) and B(53)) xor (A(109) and B(52)) xor (A(110) and B(51)) xor (A(111) and B(50)) xor (A(112) and B(49)) xor (A(113) and B(48)) xor (A(114) and B(47)) xor (A(115) and B(46)) xor (A(116) and B(45)) xor (A(117) and B(44)) xor (A(118) and B(43)) xor (A(119) and B(42)) xor (A(120) and B(41)) xor (A(121) and B(40)) xor (A(122) and B(39)) xor (A(123) and B(38)) xor (A(124) and B(37)) xor (A(125) and B(36)) xor (A(126) and B(35)) xor (A(39) and B(127)) xor (A(40) and B(126)) xor (A(41) and B(125)) xor (A(42) and B(124)) xor (A(43) and B(123)) xor (A(44) and B(122)) xor (A(45) and B(121)) xor (A(46) and B(120)) xor (A(47) and B(119)) xor (A(48) and B(118)) xor (A(49) and B(117)) xor (A(50) and B(116)) xor (A(51) and B(115)) xor (A(52) and B(114)) xor (A(53) and B(113)) xor (A(54) and B(112)) xor (A(55) and B(111)) xor (A(56) and B(110)) xor (A(57) and B(109)) xor (A(58) and B(108)) xor (A(59) and B(107)) xor (A(60) and B(106)) xor (A(61) and B(105)) xor (A(62) and B(104)) xor (A(63) and B(103)) xor (A(64) and B(102)) xor (A(65) and B(101)) xor (A(66) and B(100)) xor (A(67) and B(99)) xor (A(68) and B(98)) xor (A(69) and B(97)) xor (A(70) and B(96)) xor (A(71) and B(95)) xor (A(72) and B(94)) xor (A(73) and B(93)) xor (A(74) and B(92)) xor (A(75) and B(91)) xor (A(76) and B(90)) xor (A(77) and B(89)) xor (A(78) and B(88)) xor (A(79) and B(87)) xor (A(80) and B(86)) xor (A(81) and B(85)) xor (A(82) and B(84)) xor (A(83) and B(83)) xor (A(84) and B(82)) xor (A(85) and B(81)) xor (A(86) and B(80)) xor (A(87) and B(79)) xor (A(88) and B(78)) xor (A(89) and B(77)) xor (A(90) and B(76)) xor (A(91) and B(75)) xor (A(92) and B(74)) xor (A(93) and B(73)) xor (A(94) and B(72)) xor (A(95) and B(71)) xor (A(96) and B(70)) xor (A(97) and B(69)) xor (A(98) and B(68)) xor (A(99) and B(67)) xor (A(100) and B(66)) xor (A(101) and B(65)) xor (A(102) and B(64)) xor (A(103) and B(63)) xor (A(104) and B(62)) xor (A(105) and B(61)) xor (A(106) and B(60)) xor (A(107) and B(59)) xor (A(108) and B(58)) xor (A(109) and B(57)) xor (A(110) and B(56)) xor (A(111) and B(55)) xor (A(112) and B(54)) xor (A(113) and B(53)) xor (A(114) and B(52)) xor (A(115) and B(51)) xor (A(116) and B(50)) xor (A(117) and B(49)) xor (A(118) and B(48)) xor (A(119) and B(47)) xor (A(120) and B(46)) xor (A(121) and B(45)) xor (A(122) and B(44)) xor (A(123) and B(43)) xor (A(124) and B(42)) xor (A(125) and B(41)) xor (A(126) and B(40)) xor (A(40) and B(127)) xor (A(41) and B(126)) xor (A(42) and B(125)) xor (A(43) and B(124)) xor (A(44) and B(123)) xor (A(45) and B(122)) xor (A(46) and B(121)) xor (A(47) and B(120)) xor (A(48) and B(119)) xor (A(49) and B(118)) xor (A(50) and B(117)) xor (A(51) and B(116)) xor (A(52) and B(115)) xor (A(53) and B(114)) xor (A(54) and B(113)) xor (A(55) and B(112)) xor (A(56) and B(111)) xor (A(57) and B(110)) xor (A(58) and B(109)) xor (A(59) and B(108)) xor (A(60) and B(107)) xor (A(61) and B(106)) xor (A(62) and B(105)) xor (A(63) and B(104)) xor (A(64) and B(103)) xor (A(65) and B(102)) xor (A(66) and B(101)) xor (A(67) and B(100)) xor (A(68) and B(99)) xor (A(69) and B(98)) xor (A(70) and B(97)) xor (A(71) and B(96)) xor (A(72) and B(95)) xor (A(73) and B(94)) xor (A(74) and B(93)) xor (A(75) and B(92)) xor (A(76) and B(91)) xor (A(77) and B(90)) xor (A(78) and B(89)) xor (A(79) and B(88)) xor (A(80) and B(87)) xor (A(81) and B(86)) xor (A(82) and B(85)) xor (A(83) and B(84)) xor (A(84) and B(83)) xor (A(85) and B(82)) xor (A(86) and B(81)) xor (A(87) and B(80)) xor (A(88) and B(79)) xor (A(89) and B(78)) xor (A(90) and B(77)) xor (A(91) and B(76)) xor (A(92) and B(75)) xor (A(93) and B(74)) xor (A(94) and B(73)) xor (A(95) and B(72)) xor (A(96) and B(71)) xor (A(97) and B(70)) xor (A(98) and B(69)) xor (A(99) and B(68)) xor (A(100) and B(67)) xor (A(101) and B(66)) xor (A(102) and B(65)) xor (A(103) and B(64)) xor (A(104) and B(63)) xor (A(105) and B(62)) xor (A(106) and B(61)) xor (A(107) and B(60)) xor (A(108) and B(59)) xor (A(109) and B(58)) xor (A(110) and B(57)) xor (A(111) and B(56)) xor (A(112) and B(55)) xor (A(113) and B(54)) xor (A(114) and B(53)) xor (A(115) and B(52)) xor (A(116) and B(51)) xor (A(117) and B(50)) xor (A(118) and B(49)) xor (A(119) and B(48)) xor (A(120) and B(47)) xor (A(121) and B(46)) xor (A(122) and B(45)) xor (A(123) and B(44)) xor (A(124) and B(43)) xor (A(125) and B(42)) xor (A(126) and B(41)) xor (A(41) and B(127)) xor (A(42) and B(126)) xor (A(43) and B(125)) xor (A(44) and B(124)) xor (A(45) and B(123)) xor (A(46) and B(122)) xor (A(47) and B(121)) xor (A(48) and B(120)) xor (A(49) and B(119)) xor (A(50) and B(118)) xor (A(51) and B(117)) xor (A(52) and B(116)) xor (A(53) and B(115)) xor (A(54) and B(114)) xor (A(55) and B(113)) xor (A(56) and B(112)) xor (A(57) and B(111)) xor (A(58) and B(110)) xor (A(59) and B(109)) xor (A(60) and B(108)) xor (A(61) and B(107)) xor (A(62) and B(106)) xor (A(63) and B(105)) xor (A(64) and B(104)) xor (A(65) and B(103)) xor (A(66) and B(102)) xor (A(67) and B(101)) xor (A(68) and B(100)) xor (A(69) and B(99)) xor (A(70) and B(98)) xor (A(71) and B(97)) xor (A(72) and B(96)) xor (A(73) and B(95)) xor (A(74) and B(94)) xor (A(75) and B(93)) xor (A(76) and B(92)) xor (A(77) and B(91)) xor (A(78) and B(90)) xor (A(79) and B(89)) xor (A(80) and B(88)) xor (A(81) and B(87)) xor (A(82) and B(86)) xor (A(83) and B(85)) xor (A(84) and B(84)) xor (A(85) and B(83)) xor (A(86) and B(82)) xor (A(87) and B(81)) xor (A(88) and B(80)) xor (A(89) and B(79)) xor (A(90) and B(78)) xor (A(91) and B(77)) xor (A(92) and B(76)) xor (A(93) and B(75)) xor (A(94) and B(74)) xor (A(95) and B(73)) xor (A(96) and B(72)) xor (A(97) and B(71)) xor (A(98) and B(70)) xor (A(99) and B(69)) xor (A(100) and B(68)) xor (A(101) and B(67)) xor (A(102) and B(66)) xor (A(103) and B(65)) xor (A(104) and B(64)) xor (A(105) and B(63)) xor (A(106) and B(62)) xor (A(107) and B(61)) xor (A(108) and B(60)) xor (A(109) and B(59)) xor (A(110) and B(58)) xor (A(111) and B(57)) xor (A(112) and B(56)) xor (A(113) and B(55)) xor (A(114) and B(54)) xor (A(115) and B(53)) xor (A(116) and B(52)) xor (A(117) and B(51)) xor (A(118) and B(50)) xor (A(119) and B(49)) xor (A(120) and B(48)) xor (A(121) and B(47)) xor (A(122) and B(46)) xor (A(123) and B(45)) xor (A(124) and B(44)) xor (A(125) and B(43)) xor (A(126) and B(43));
    C(42)  <= (A(0) and B(42)) xor (A(1) and B(41)) xor (A(2) and B(40)) xor (A(3) and B(39)) xor (A(4) and B(38)) xor (A(5) and B(37)) xor (A(6) and B(36)) xor (A(7) and B(35)) xor (A(8) and B(34)) xor (A(9) and B(33)) xor (A(10) and B(32)) xor (A(11) and B(31)) xor (A(12) and B(30)) xor (A(13) and B(29)) xor (A(14) and B(28)) xor (A(15) and B(27)) xor (A(16) and B(26)) xor (A(17) and B(25)) xor (A(18) and B(24)) xor (A(19) and B(23)) xor (A(20) and B(23)) xor (A(21) and B(21)) xor (A(23) and B(20)) xor (A(23) and B(19)) xor (A(24) and B(18)) xor (A(25) and B(17)) xor (A(26) and B(16)) xor (A(27) and B(15)) xor (A(28) and B(14)) xor (A(29) and B(13)) xor (A(30) and B(12)) xor (A(31) and B(11)) xor (A(32) and B(10)) xor (A(33) and B(9)) xor (A(34) and B(8)) xor (A(35) and B(7)) xor (A(36) and B(6)) xor (A(37) and B(5)) xor (A(38) and B(4)) xor (A(39) and B(3)) xor (A(40) and B(2)) xor (A(41) and B(1)) xor (A(42) and B(0)) xor (A(35) and B(127)) xor (A(36) and B(126)) xor (A(37) and B(125)) xor (A(38) and B(124)) xor (A(39) and B(123)) xor (A(40) and B(122)) xor (A(41) and B(121)) xor (A(42) and B(120)) xor (A(43) and B(119)) xor (A(44) and B(118)) xor (A(45) and B(117)) xor (A(46) and B(116)) xor (A(47) and B(115)) xor (A(48) and B(114)) xor (A(49) and B(113)) xor (A(50) and B(112)) xor (A(51) and B(111)) xor (A(52) and B(110)) xor (A(53) and B(109)) xor (A(54) and B(108)) xor (A(55) and B(107)) xor (A(56) and B(106)) xor (A(57) and B(105)) xor (A(58) and B(104)) xor (A(59) and B(103)) xor (A(60) and B(102)) xor (A(61) and B(101)) xor (A(62) and B(100)) xor (A(63) and B(99)) xor (A(64) and B(98)) xor (A(65) and B(97)) xor (A(66) and B(96)) xor (A(67) and B(95)) xor (A(68) and B(94)) xor (A(69) and B(93)) xor (A(70) and B(92)) xor (A(71) and B(91)) xor (A(72) and B(90)) xor (A(73) and B(89)) xor (A(74) and B(88)) xor (A(75) and B(87)) xor (A(76) and B(86)) xor (A(77) and B(85)) xor (A(78) and B(84)) xor (A(79) and B(83)) xor (A(80) and B(82)) xor (A(81) and B(81)) xor (A(82) and B(80)) xor (A(83) and B(79)) xor (A(84) and B(78)) xor (A(85) and B(77)) xor (A(86) and B(76)) xor (A(87) and B(75)) xor (A(88) and B(74)) xor (A(89) and B(73)) xor (A(90) and B(72)) xor (A(91) and B(71)) xor (A(92) and B(70)) xor (A(93) and B(69)) xor (A(94) and B(68)) xor (A(95) and B(67)) xor (A(96) and B(66)) xor (A(97) and B(65)) xor (A(98) and B(64)) xor (A(99) and B(63)) xor (A(100) and B(62)) xor (A(101) and B(61)) xor (A(102) and B(60)) xor (A(103) and B(59)) xor (A(104) and B(58)) xor (A(105) and B(57)) xor (A(106) and B(56)) xor (A(107) and B(55)) xor (A(108) and B(54)) xor (A(109) and B(53)) xor (A(110) and B(52)) xor (A(111) and B(51)) xor (A(112) and B(50)) xor (A(113) and B(49)) xor (A(114) and B(48)) xor (A(115) and B(47)) xor (A(116) and B(46)) xor (A(117) and B(45)) xor (A(118) and B(44)) xor (A(119) and B(43)) xor (A(120) and B(42)) xor (A(121) and B(41)) xor (A(122) and B(40)) xor (A(123) and B(39)) xor (A(124) and B(38)) xor (A(125) and B(37)) xor (A(126) and B(36)) xor (A(40) and B(127)) xor (A(41) and B(126)) xor (A(42) and B(125)) xor (A(43) and B(124)) xor (A(44) and B(123)) xor (A(45) and B(122)) xor (A(46) and B(121)) xor (A(47) and B(120)) xor (A(48) and B(119)) xor (A(49) and B(118)) xor (A(50) and B(117)) xor (A(51) and B(116)) xor (A(52) and B(115)) xor (A(53) and B(114)) xor (A(54) and B(113)) xor (A(55) and B(112)) xor (A(56) and B(111)) xor (A(57) and B(110)) xor (A(58) and B(109)) xor (A(59) and B(108)) xor (A(60) and B(107)) xor (A(61) and B(106)) xor (A(62) and B(105)) xor (A(63) and B(104)) xor (A(64) and B(103)) xor (A(65) and B(102)) xor (A(66) and B(101)) xor (A(67) and B(100)) xor (A(68) and B(99)) xor (A(69) and B(98)) xor (A(70) and B(97)) xor (A(71) and B(96)) xor (A(72) and B(95)) xor (A(73) and B(94)) xor (A(74) and B(93)) xor (A(75) and B(92)) xor (A(76) and B(91)) xor (A(77) and B(90)) xor (A(78) and B(89)) xor (A(79) and B(88)) xor (A(80) and B(87)) xor (A(81) and B(86)) xor (A(82) and B(85)) xor (A(83) and B(84)) xor (A(84) and B(83)) xor (A(85) and B(82)) xor (A(86) and B(81)) xor (A(87) and B(80)) xor (A(88) and B(79)) xor (A(89) and B(78)) xor (A(90) and B(77)) xor (A(91) and B(76)) xor (A(92) and B(75)) xor (A(93) and B(74)) xor (A(94) and B(73)) xor (A(95) and B(72)) xor (A(96) and B(71)) xor (A(97) and B(70)) xor (A(98) and B(69)) xor (A(99) and B(68)) xor (A(100) and B(67)) xor (A(101) and B(66)) xor (A(102) and B(65)) xor (A(103) and B(64)) xor (A(104) and B(63)) xor (A(105) and B(62)) xor (A(106) and B(61)) xor (A(107) and B(60)) xor (A(108) and B(59)) xor (A(109) and B(58)) xor (A(110) and B(57)) xor (A(111) and B(56)) xor (A(112) and B(55)) xor (A(113) and B(54)) xor (A(114) and B(53)) xor (A(115) and B(52)) xor (A(116) and B(51)) xor (A(117) and B(50)) xor (A(118) and B(49)) xor (A(119) and B(48)) xor (A(120) and B(47)) xor (A(121) and B(46)) xor (A(122) and B(45)) xor (A(123) and B(44)) xor (A(124) and B(43)) xor (A(125) and B(42)) xor (A(126) and B(41)) xor (A(41) and B(127)) xor (A(42) and B(126)) xor (A(43) and B(125)) xor (A(44) and B(124)) xor (A(45) and B(123)) xor (A(46) and B(122)) xor (A(47) and B(121)) xor (A(48) and B(120)) xor (A(49) and B(119)) xor (A(50) and B(118)) xor (A(51) and B(117)) xor (A(52) and B(116)) xor (A(53) and B(115)) xor (A(54) and B(114)) xor (A(55) and B(113)) xor (A(56) and B(112)) xor (A(57) and B(111)) xor (A(58) and B(110)) xor (A(59) and B(109)) xor (A(60) and B(108)) xor (A(61) and B(107)) xor (A(62) and B(106)) xor (A(63) and B(105)) xor (A(64) and B(104)) xor (A(65) and B(103)) xor (A(66) and B(102)) xor (A(67) and B(101)) xor (A(68) and B(100)) xor (A(69) and B(99)) xor (A(70) and B(98)) xor (A(71) and B(97)) xor (A(72) and B(96)) xor (A(73) and B(95)) xor (A(74) and B(94)) xor (A(75) and B(93)) xor (A(76) and B(92)) xor (A(77) and B(91)) xor (A(78) and B(90)) xor (A(79) and B(89)) xor (A(80) and B(88)) xor (A(81) and B(87)) xor (A(82) and B(86)) xor (A(83) and B(85)) xor (A(84) and B(84)) xor (A(85) and B(83)) xor (A(86) and B(82)) xor (A(87) and B(81)) xor (A(88) and B(80)) xor (A(89) and B(79)) xor (A(90) and B(78)) xor (A(91) and B(77)) xor (A(92) and B(76)) xor (A(93) and B(75)) xor (A(94) and B(74)) xor (A(95) and B(73)) xor (A(96) and B(72)) xor (A(97) and B(71)) xor (A(98) and B(70)) xor (A(99) and B(69)) xor (A(100) and B(68)) xor (A(101) and B(67)) xor (A(102) and B(66)) xor (A(103) and B(65)) xor (A(104) and B(64)) xor (A(105) and B(63)) xor (A(106) and B(62)) xor (A(107) and B(61)) xor (A(108) and B(60)) xor (A(109) and B(59)) xor (A(110) and B(58)) xor (A(111) and B(57)) xor (A(112) and B(56)) xor (A(113) and B(55)) xor (A(114) and B(54)) xor (A(115) and B(53)) xor (A(116) and B(52)) xor (A(117) and B(51)) xor (A(118) and B(50)) xor (A(119) and B(49)) xor (A(120) and B(48)) xor (A(121) and B(47)) xor (A(122) and B(46)) xor (A(123) and B(45)) xor (A(124) and B(44)) xor (A(125) and B(43)) xor (A(126) and B(42)) xor (A(42) and B(127)) xor (A(43) and B(126)) xor (A(44) and B(125)) xor (A(45) and B(124)) xor (A(46) and B(123)) xor (A(47) and B(122)) xor (A(48) and B(121)) xor (A(49) and B(120)) xor (A(50) and B(119)) xor (A(51) and B(118)) xor (A(52) and B(117)) xor (A(53) and B(116)) xor (A(54) and B(115)) xor (A(55) and B(114)) xor (A(56) and B(113)) xor (A(57) and B(112)) xor (A(58) and B(111)) xor (A(59) and B(110)) xor (A(60) and B(109)) xor (A(61) and B(108)) xor (A(62) and B(107)) xor (A(63) and B(106)) xor (A(64) and B(105)) xor (A(65) and B(104)) xor (A(66) and B(103)) xor (A(67) and B(102)) xor (A(68) and B(101)) xor (A(69) and B(100)) xor (A(70) and B(99)) xor (A(71) and B(98)) xor (A(72) and B(97)) xor (A(73) and B(96)) xor (A(74) and B(95)) xor (A(75) and B(94)) xor (A(76) and B(93)) xor (A(77) and B(92)) xor (A(78) and B(91)) xor (A(79) and B(90)) xor (A(80) and B(89)) xor (A(81) and B(88)) xor (A(82) and B(87)) xor (A(83) and B(86)) xor (A(84) and B(85)) xor (A(85) and B(84)) xor (A(86) and B(83)) xor (A(87) and B(82)) xor (A(88) and B(81)) xor (A(89) and B(80)) xor (A(90) and B(79)) xor (A(91) and B(78)) xor (A(92) and B(77)) xor (A(93) and B(76)) xor (A(94) and B(75)) xor (A(95) and B(74)) xor (A(96) and B(73)) xor (A(97) and B(72)) xor (A(98) and B(71)) xor (A(99) and B(70)) xor (A(100) and B(69)) xor (A(101) and B(68)) xor (A(102) and B(67)) xor (A(103) and B(66)) xor (A(104) and B(65)) xor (A(105) and B(64)) xor (A(106) and B(63)) xor (A(107) and B(62)) xor (A(108) and B(61)) xor (A(109) and B(60)) xor (A(110) and B(59)) xor (A(111) and B(58)) xor (A(112) and B(57)) xor (A(113) and B(56)) xor (A(114) and B(55)) xor (A(115) and B(54)) xor (A(116) and B(53)) xor (A(117) and B(52)) xor (A(118) and B(51)) xor (A(119) and B(50)) xor (A(120) and B(49)) xor (A(121) and B(48)) xor (A(122) and B(47)) xor (A(123) and B(46)) xor (A(124) and B(45)) xor (A(125) and B(44)) xor (A(126) and B(44));
    C(43)  <= (A(0) and B(43)) xor (A(1) and B(42)) xor (A(2) and B(41)) xor (A(3) and B(40)) xor (A(4) and B(39)) xor (A(5) and B(38)) xor (A(6) and B(37)) xor (A(7) and B(36)) xor (A(8) and B(35)) xor (A(9) and B(34)) xor (A(10) and B(33)) xor (A(11) and B(32)) xor (A(12) and B(31)) xor (A(13) and B(30)) xor (A(14) and B(29)) xor (A(15) and B(28)) xor (A(16) and B(27)) xor (A(17) and B(26)) xor (A(18) and B(25)) xor (A(19) and B(24)) xor (A(20) and B(23)) xor (A(21) and B(23)) xor (A(23) and B(21)) xor (A(23) and B(20)) xor (A(24) and B(19)) xor (A(25) and B(18)) xor (A(26) and B(17)) xor (A(27) and B(16)) xor (A(28) and B(15)) xor (A(29) and B(14)) xor (A(30) and B(13)) xor (A(31) and B(12)) xor (A(32) and B(11)) xor (A(33) and B(10)) xor (A(34) and B(9)) xor (A(35) and B(8)) xor (A(36) and B(7)) xor (A(37) and B(6)) xor (A(38) and B(5)) xor (A(39) and B(4)) xor (A(40) and B(3)) xor (A(41) and B(2)) xor (A(42) and B(1)) xor (A(43) and B(0)) xor (A(36) and B(127)) xor (A(37) and B(126)) xor (A(38) and B(125)) xor (A(39) and B(124)) xor (A(40) and B(123)) xor (A(41) and B(122)) xor (A(42) and B(121)) xor (A(43) and B(120)) xor (A(44) and B(119)) xor (A(45) and B(118)) xor (A(46) and B(117)) xor (A(47) and B(116)) xor (A(48) and B(115)) xor (A(49) and B(114)) xor (A(50) and B(113)) xor (A(51) and B(112)) xor (A(52) and B(111)) xor (A(53) and B(110)) xor (A(54) and B(109)) xor (A(55) and B(108)) xor (A(56) and B(107)) xor (A(57) and B(106)) xor (A(58) and B(105)) xor (A(59) and B(104)) xor (A(60) and B(103)) xor (A(61) and B(102)) xor (A(62) and B(101)) xor (A(63) and B(100)) xor (A(64) and B(99)) xor (A(65) and B(98)) xor (A(66) and B(97)) xor (A(67) and B(96)) xor (A(68) and B(95)) xor (A(69) and B(94)) xor (A(70) and B(93)) xor (A(71) and B(92)) xor (A(72) and B(91)) xor (A(73) and B(90)) xor (A(74) and B(89)) xor (A(75) and B(88)) xor (A(76) and B(87)) xor (A(77) and B(86)) xor (A(78) and B(85)) xor (A(79) and B(84)) xor (A(80) and B(83)) xor (A(81) and B(82)) xor (A(82) and B(81)) xor (A(83) and B(80)) xor (A(84) and B(79)) xor (A(85) and B(78)) xor (A(86) and B(77)) xor (A(87) and B(76)) xor (A(88) and B(75)) xor (A(89) and B(74)) xor (A(90) and B(73)) xor (A(91) and B(72)) xor (A(92) and B(71)) xor (A(93) and B(70)) xor (A(94) and B(69)) xor (A(95) and B(68)) xor (A(96) and B(67)) xor (A(97) and B(66)) xor (A(98) and B(65)) xor (A(99) and B(64)) xor (A(100) and B(63)) xor (A(101) and B(62)) xor (A(102) and B(61)) xor (A(103) and B(60)) xor (A(104) and B(59)) xor (A(105) and B(58)) xor (A(106) and B(57)) xor (A(107) and B(56)) xor (A(108) and B(55)) xor (A(109) and B(54)) xor (A(110) and B(53)) xor (A(111) and B(52)) xor (A(112) and B(51)) xor (A(113) and B(50)) xor (A(114) and B(49)) xor (A(115) and B(48)) xor (A(116) and B(47)) xor (A(117) and B(46)) xor (A(118) and B(45)) xor (A(119) and B(44)) xor (A(120) and B(43)) xor (A(121) and B(42)) xor (A(122) and B(41)) xor (A(123) and B(40)) xor (A(124) and B(39)) xor (A(125) and B(38)) xor (A(126) and B(37)) xor (A(41) and B(127)) xor (A(42) and B(126)) xor (A(43) and B(125)) xor (A(44) and B(124)) xor (A(45) and B(123)) xor (A(46) and B(122)) xor (A(47) and B(121)) xor (A(48) and B(120)) xor (A(49) and B(119)) xor (A(50) and B(118)) xor (A(51) and B(117)) xor (A(52) and B(116)) xor (A(53) and B(115)) xor (A(54) and B(114)) xor (A(55) and B(113)) xor (A(56) and B(112)) xor (A(57) and B(111)) xor (A(58) and B(110)) xor (A(59) and B(109)) xor (A(60) and B(108)) xor (A(61) and B(107)) xor (A(62) and B(106)) xor (A(63) and B(105)) xor (A(64) and B(104)) xor (A(65) and B(103)) xor (A(66) and B(102)) xor (A(67) and B(101)) xor (A(68) and B(100)) xor (A(69) and B(99)) xor (A(70) and B(98)) xor (A(71) and B(97)) xor (A(72) and B(96)) xor (A(73) and B(95)) xor (A(74) and B(94)) xor (A(75) and B(93)) xor (A(76) and B(92)) xor (A(77) and B(91)) xor (A(78) and B(90)) xor (A(79) and B(89)) xor (A(80) and B(88)) xor (A(81) and B(87)) xor (A(82) and B(86)) xor (A(83) and B(85)) xor (A(84) and B(84)) xor (A(85) and B(83)) xor (A(86) and B(82)) xor (A(87) and B(81)) xor (A(88) and B(80)) xor (A(89) and B(79)) xor (A(90) and B(78)) xor (A(91) and B(77)) xor (A(92) and B(76)) xor (A(93) and B(75)) xor (A(94) and B(74)) xor (A(95) and B(73)) xor (A(96) and B(72)) xor (A(97) and B(71)) xor (A(98) and B(70)) xor (A(99) and B(69)) xor (A(100) and B(68)) xor (A(101) and B(67)) xor (A(102) and B(66)) xor (A(103) and B(65)) xor (A(104) and B(64)) xor (A(105) and B(63)) xor (A(106) and B(62)) xor (A(107) and B(61)) xor (A(108) and B(60)) xor (A(109) and B(59)) xor (A(110) and B(58)) xor (A(111) and B(57)) xor (A(112) and B(56)) xor (A(113) and B(55)) xor (A(114) and B(54)) xor (A(115) and B(53)) xor (A(116) and B(52)) xor (A(117) and B(51)) xor (A(118) and B(50)) xor (A(119) and B(49)) xor (A(120) and B(48)) xor (A(121) and B(47)) xor (A(122) and B(46)) xor (A(123) and B(45)) xor (A(124) and B(44)) xor (A(125) and B(43)) xor (A(126) and B(42)) xor (A(42) and B(127)) xor (A(43) and B(126)) xor (A(44) and B(125)) xor (A(45) and B(124)) xor (A(46) and B(123)) xor (A(47) and B(122)) xor (A(48) and B(121)) xor (A(49) and B(120)) xor (A(50) and B(119)) xor (A(51) and B(118)) xor (A(52) and B(117)) xor (A(53) and B(116)) xor (A(54) and B(115)) xor (A(55) and B(114)) xor (A(56) and B(113)) xor (A(57) and B(112)) xor (A(58) and B(111)) xor (A(59) and B(110)) xor (A(60) and B(109)) xor (A(61) and B(108)) xor (A(62) and B(107)) xor (A(63) and B(106)) xor (A(64) and B(105)) xor (A(65) and B(104)) xor (A(66) and B(103)) xor (A(67) and B(102)) xor (A(68) and B(101)) xor (A(69) and B(100)) xor (A(70) and B(99)) xor (A(71) and B(98)) xor (A(72) and B(97)) xor (A(73) and B(96)) xor (A(74) and B(95)) xor (A(75) and B(94)) xor (A(76) and B(93)) xor (A(77) and B(92)) xor (A(78) and B(91)) xor (A(79) and B(90)) xor (A(80) and B(89)) xor (A(81) and B(88)) xor (A(82) and B(87)) xor (A(83) and B(86)) xor (A(84) and B(85)) xor (A(85) and B(84)) xor (A(86) and B(83)) xor (A(87) and B(82)) xor (A(88) and B(81)) xor (A(89) and B(80)) xor (A(90) and B(79)) xor (A(91) and B(78)) xor (A(92) and B(77)) xor (A(93) and B(76)) xor (A(94) and B(75)) xor (A(95) and B(74)) xor (A(96) and B(73)) xor (A(97) and B(72)) xor (A(98) and B(71)) xor (A(99) and B(70)) xor (A(100) and B(69)) xor (A(101) and B(68)) xor (A(102) and B(67)) xor (A(103) and B(66)) xor (A(104) and B(65)) xor (A(105) and B(64)) xor (A(106) and B(63)) xor (A(107) and B(62)) xor (A(108) and B(61)) xor (A(109) and B(60)) xor (A(110) and B(59)) xor (A(111) and B(58)) xor (A(112) and B(57)) xor (A(113) and B(56)) xor (A(114) and B(55)) xor (A(115) and B(54)) xor (A(116) and B(53)) xor (A(117) and B(52)) xor (A(118) and B(51)) xor (A(119) and B(50)) xor (A(120) and B(49)) xor (A(121) and B(48)) xor (A(122) and B(47)) xor (A(123) and B(46)) xor (A(124) and B(45)) xor (A(125) and B(44)) xor (A(126) and B(43)) xor (A(43) and B(127)) xor (A(44) and B(126)) xor (A(45) and B(125)) xor (A(46) and B(124)) xor (A(47) and B(123)) xor (A(48) and B(122)) xor (A(49) and B(121)) xor (A(50) and B(120)) xor (A(51) and B(119)) xor (A(52) and B(118)) xor (A(53) and B(117)) xor (A(54) and B(116)) xor (A(55) and B(115)) xor (A(56) and B(114)) xor (A(57) and B(113)) xor (A(58) and B(112)) xor (A(59) and B(111)) xor (A(60) and B(110)) xor (A(61) and B(109)) xor (A(62) and B(108)) xor (A(63) and B(107)) xor (A(64) and B(106)) xor (A(65) and B(105)) xor (A(66) and B(104)) xor (A(67) and B(103)) xor (A(68) and B(102)) xor (A(69) and B(101)) xor (A(70) and B(100)) xor (A(71) and B(99)) xor (A(72) and B(98)) xor (A(73) and B(97)) xor (A(74) and B(96)) xor (A(75) and B(95)) xor (A(76) and B(94)) xor (A(77) and B(93)) xor (A(78) and B(92)) xor (A(79) and B(91)) xor (A(80) and B(90)) xor (A(81) and B(89)) xor (A(82) and B(88)) xor (A(83) and B(87)) xor (A(84) and B(86)) xor (A(85) and B(85)) xor (A(86) and B(84)) xor (A(87) and B(83)) xor (A(88) and B(82)) xor (A(89) and B(81)) xor (A(90) and B(80)) xor (A(91) and B(79)) xor (A(92) and B(78)) xor (A(93) and B(77)) xor (A(94) and B(76)) xor (A(95) and B(75)) xor (A(96) and B(74)) xor (A(97) and B(73)) xor (A(98) and B(72)) xor (A(99) and B(71)) xor (A(100) and B(70)) xor (A(101) and B(69)) xor (A(102) and B(68)) xor (A(103) and B(67)) xor (A(104) and B(66)) xor (A(105) and B(65)) xor (A(106) and B(64)) xor (A(107) and B(63)) xor (A(108) and B(62)) xor (A(109) and B(61)) xor (A(110) and B(60)) xor (A(111) and B(59)) xor (A(112) and B(58)) xor (A(113) and B(57)) xor (A(114) and B(56)) xor (A(115) and B(55)) xor (A(116) and B(54)) xor (A(117) and B(53)) xor (A(118) and B(52)) xor (A(119) and B(51)) xor (A(120) and B(50)) xor (A(121) and B(49)) xor (A(122) and B(48)) xor (A(123) and B(47)) xor (A(124) and B(46)) xor (A(125) and B(45)) xor (A(126) and B(45));
    C(44)  <= (A(0) and B(44)) xor (A(1) and B(43)) xor (A(2) and B(42)) xor (A(3) and B(41)) xor (A(4) and B(40)) xor (A(5) and B(39)) xor (A(6) and B(38)) xor (A(7) and B(37)) xor (A(8) and B(36)) xor (A(9) and B(35)) xor (A(10) and B(34)) xor (A(11) and B(33)) xor (A(12) and B(32)) xor (A(13) and B(31)) xor (A(14) and B(30)) xor (A(15) and B(29)) xor (A(16) and B(28)) xor (A(17) and B(27)) xor (A(18) and B(26)) xor (A(19) and B(25)) xor (A(20) and B(24)) xor (A(21) and B(23)) xor (A(23) and B(23)) xor (A(23) and B(21)) xor (A(24) and B(20)) xor (A(25) and B(19)) xor (A(26) and B(18)) xor (A(27) and B(17)) xor (A(28) and B(16)) xor (A(29) and B(15)) xor (A(30) and B(14)) xor (A(31) and B(13)) xor (A(32) and B(12)) xor (A(33) and B(11)) xor (A(34) and B(10)) xor (A(35) and B(9)) xor (A(36) and B(8)) xor (A(37) and B(7)) xor (A(38) and B(6)) xor (A(39) and B(5)) xor (A(40) and B(4)) xor (A(41) and B(3)) xor (A(42) and B(2)) xor (A(43) and B(1)) xor (A(44) and B(0)) xor (A(37) and B(127)) xor (A(38) and B(126)) xor (A(39) and B(125)) xor (A(40) and B(124)) xor (A(41) and B(123)) xor (A(42) and B(122)) xor (A(43) and B(121)) xor (A(44) and B(120)) xor (A(45) and B(119)) xor (A(46) and B(118)) xor (A(47) and B(117)) xor (A(48) and B(116)) xor (A(49) and B(115)) xor (A(50) and B(114)) xor (A(51) and B(113)) xor (A(52) and B(112)) xor (A(53) and B(111)) xor (A(54) and B(110)) xor (A(55) and B(109)) xor (A(56) and B(108)) xor (A(57) and B(107)) xor (A(58) and B(106)) xor (A(59) and B(105)) xor (A(60) and B(104)) xor (A(61) and B(103)) xor (A(62) and B(102)) xor (A(63) and B(101)) xor (A(64) and B(100)) xor (A(65) and B(99)) xor (A(66) and B(98)) xor (A(67) and B(97)) xor (A(68) and B(96)) xor (A(69) and B(95)) xor (A(70) and B(94)) xor (A(71) and B(93)) xor (A(72) and B(92)) xor (A(73) and B(91)) xor (A(74) and B(90)) xor (A(75) and B(89)) xor (A(76) and B(88)) xor (A(77) and B(87)) xor (A(78) and B(86)) xor (A(79) and B(85)) xor (A(80) and B(84)) xor (A(81) and B(83)) xor (A(82) and B(82)) xor (A(83) and B(81)) xor (A(84) and B(80)) xor (A(85) and B(79)) xor (A(86) and B(78)) xor (A(87) and B(77)) xor (A(88) and B(76)) xor (A(89) and B(75)) xor (A(90) and B(74)) xor (A(91) and B(73)) xor (A(92) and B(72)) xor (A(93) and B(71)) xor (A(94) and B(70)) xor (A(95) and B(69)) xor (A(96) and B(68)) xor (A(97) and B(67)) xor (A(98) and B(66)) xor (A(99) and B(65)) xor (A(100) and B(64)) xor (A(101) and B(63)) xor (A(102) and B(62)) xor (A(103) and B(61)) xor (A(104) and B(60)) xor (A(105) and B(59)) xor (A(106) and B(58)) xor (A(107) and B(57)) xor (A(108) and B(56)) xor (A(109) and B(55)) xor (A(110) and B(54)) xor (A(111) and B(53)) xor (A(112) and B(52)) xor (A(113) and B(51)) xor (A(114) and B(50)) xor (A(115) and B(49)) xor (A(116) and B(48)) xor (A(117) and B(47)) xor (A(118) and B(46)) xor (A(119) and B(45)) xor (A(120) and B(44)) xor (A(121) and B(43)) xor (A(122) and B(42)) xor (A(123) and B(41)) xor (A(124) and B(40)) xor (A(125) and B(39)) xor (A(126) and B(38)) xor (A(42) and B(127)) xor (A(43) and B(126)) xor (A(44) and B(125)) xor (A(45) and B(124)) xor (A(46) and B(123)) xor (A(47) and B(122)) xor (A(48) and B(121)) xor (A(49) and B(120)) xor (A(50) and B(119)) xor (A(51) and B(118)) xor (A(52) and B(117)) xor (A(53) and B(116)) xor (A(54) and B(115)) xor (A(55) and B(114)) xor (A(56) and B(113)) xor (A(57) and B(112)) xor (A(58) and B(111)) xor (A(59) and B(110)) xor (A(60) and B(109)) xor (A(61) and B(108)) xor (A(62) and B(107)) xor (A(63) and B(106)) xor (A(64) and B(105)) xor (A(65) and B(104)) xor (A(66) and B(103)) xor (A(67) and B(102)) xor (A(68) and B(101)) xor (A(69) and B(100)) xor (A(70) and B(99)) xor (A(71) and B(98)) xor (A(72) and B(97)) xor (A(73) and B(96)) xor (A(74) and B(95)) xor (A(75) and B(94)) xor (A(76) and B(93)) xor (A(77) and B(92)) xor (A(78) and B(91)) xor (A(79) and B(90)) xor (A(80) and B(89)) xor (A(81) and B(88)) xor (A(82) and B(87)) xor (A(83) and B(86)) xor (A(84) and B(85)) xor (A(85) and B(84)) xor (A(86) and B(83)) xor (A(87) and B(82)) xor (A(88) and B(81)) xor (A(89) and B(80)) xor (A(90) and B(79)) xor (A(91) and B(78)) xor (A(92) and B(77)) xor (A(93) and B(76)) xor (A(94) and B(75)) xor (A(95) and B(74)) xor (A(96) and B(73)) xor (A(97) and B(72)) xor (A(98) and B(71)) xor (A(99) and B(70)) xor (A(100) and B(69)) xor (A(101) and B(68)) xor (A(102) and B(67)) xor (A(103) and B(66)) xor (A(104) and B(65)) xor (A(105) and B(64)) xor (A(106) and B(63)) xor (A(107) and B(62)) xor (A(108) and B(61)) xor (A(109) and B(60)) xor (A(110) and B(59)) xor (A(111) and B(58)) xor (A(112) and B(57)) xor (A(113) and B(56)) xor (A(114) and B(55)) xor (A(115) and B(54)) xor (A(116) and B(53)) xor (A(117) and B(52)) xor (A(118) and B(51)) xor (A(119) and B(50)) xor (A(120) and B(49)) xor (A(121) and B(48)) xor (A(122) and B(47)) xor (A(123) and B(46)) xor (A(124) and B(45)) xor (A(125) and B(44)) xor (A(126) and B(43)) xor (A(43) and B(127)) xor (A(44) and B(126)) xor (A(45) and B(125)) xor (A(46) and B(124)) xor (A(47) and B(123)) xor (A(48) and B(122)) xor (A(49) and B(121)) xor (A(50) and B(120)) xor (A(51) and B(119)) xor (A(52) and B(118)) xor (A(53) and B(117)) xor (A(54) and B(116)) xor (A(55) and B(115)) xor (A(56) and B(114)) xor (A(57) and B(113)) xor (A(58) and B(112)) xor (A(59) and B(111)) xor (A(60) and B(110)) xor (A(61) and B(109)) xor (A(62) and B(108)) xor (A(63) and B(107)) xor (A(64) and B(106)) xor (A(65) and B(105)) xor (A(66) and B(104)) xor (A(67) and B(103)) xor (A(68) and B(102)) xor (A(69) and B(101)) xor (A(70) and B(100)) xor (A(71) and B(99)) xor (A(72) and B(98)) xor (A(73) and B(97)) xor (A(74) and B(96)) xor (A(75) and B(95)) xor (A(76) and B(94)) xor (A(77) and B(93)) xor (A(78) and B(92)) xor (A(79) and B(91)) xor (A(80) and B(90)) xor (A(81) and B(89)) xor (A(82) and B(88)) xor (A(83) and B(87)) xor (A(84) and B(86)) xor (A(85) and B(85)) xor (A(86) and B(84)) xor (A(87) and B(83)) xor (A(88) and B(82)) xor (A(89) and B(81)) xor (A(90) and B(80)) xor (A(91) and B(79)) xor (A(92) and B(78)) xor (A(93) and B(77)) xor (A(94) and B(76)) xor (A(95) and B(75)) xor (A(96) and B(74)) xor (A(97) and B(73)) xor (A(98) and B(72)) xor (A(99) and B(71)) xor (A(100) and B(70)) xor (A(101) and B(69)) xor (A(102) and B(68)) xor (A(103) and B(67)) xor (A(104) and B(66)) xor (A(105) and B(65)) xor (A(106) and B(64)) xor (A(107) and B(63)) xor (A(108) and B(62)) xor (A(109) and B(61)) xor (A(110) and B(60)) xor (A(111) and B(59)) xor (A(112) and B(58)) xor (A(113) and B(57)) xor (A(114) and B(56)) xor (A(115) and B(55)) xor (A(116) and B(54)) xor (A(117) and B(53)) xor (A(118) and B(52)) xor (A(119) and B(51)) xor (A(120) and B(50)) xor (A(121) and B(49)) xor (A(122) and B(48)) xor (A(123) and B(47)) xor (A(124) and B(46)) xor (A(125) and B(45)) xor (A(126) and B(44)) xor (A(44) and B(127)) xor (A(45) and B(126)) xor (A(46) and B(125)) xor (A(47) and B(124)) xor (A(48) and B(123)) xor (A(49) and B(122)) xor (A(50) and B(121)) xor (A(51) and B(120)) xor (A(52) and B(119)) xor (A(53) and B(118)) xor (A(54) and B(117)) xor (A(55) and B(116)) xor (A(56) and B(115)) xor (A(57) and B(114)) xor (A(58) and B(113)) xor (A(59) and B(112)) xor (A(60) and B(111)) xor (A(61) and B(110)) xor (A(62) and B(109)) xor (A(63) and B(108)) xor (A(64) and B(107)) xor (A(65) and B(106)) xor (A(66) and B(105)) xor (A(67) and B(104)) xor (A(68) and B(103)) xor (A(69) and B(102)) xor (A(70) and B(101)) xor (A(71) and B(100)) xor (A(72) and B(99)) xor (A(73) and B(98)) xor (A(74) and B(97)) xor (A(75) and B(96)) xor (A(76) and B(95)) xor (A(77) and B(94)) xor (A(78) and B(93)) xor (A(79) and B(92)) xor (A(80) and B(91)) xor (A(81) and B(90)) xor (A(82) and B(89)) xor (A(83) and B(88)) xor (A(84) and B(87)) xor (A(85) and B(86)) xor (A(86) and B(85)) xor (A(87) and B(84)) xor (A(88) and B(83)) xor (A(89) and B(82)) xor (A(90) and B(81)) xor (A(91) and B(80)) xor (A(92) and B(79)) xor (A(93) and B(78)) xor (A(94) and B(77)) xor (A(95) and B(76)) xor (A(96) and B(75)) xor (A(97) and B(74)) xor (A(98) and B(73)) xor (A(99) and B(72)) xor (A(100) and B(71)) xor (A(101) and B(70)) xor (A(102) and B(69)) xor (A(103) and B(68)) xor (A(104) and B(67)) xor (A(105) and B(66)) xor (A(106) and B(65)) xor (A(107) and B(64)) xor (A(108) and B(63)) xor (A(109) and B(62)) xor (A(110) and B(61)) xor (A(111) and B(60)) xor (A(112) and B(59)) xor (A(113) and B(58)) xor (A(114) and B(57)) xor (A(115) and B(56)) xor (A(116) and B(55)) xor (A(117) and B(54)) xor (A(118) and B(53)) xor (A(119) and B(52)) xor (A(120) and B(51)) xor (A(121) and B(50)) xor (A(122) and B(49)) xor (A(123) and B(48)) xor (A(124) and B(47)) xor (A(125) and B(46)) xor (A(126) and B(46));
    C(45)  <= (A(0) and B(45)) xor (A(1) and B(44)) xor (A(2) and B(43)) xor (A(3) and B(42)) xor (A(4) and B(41)) xor (A(5) and B(40)) xor (A(6) and B(39)) xor (A(7) and B(38)) xor (A(8) and B(37)) xor (A(9) and B(36)) xor (A(10) and B(35)) xor (A(11) and B(34)) xor (A(12) and B(33)) xor (A(13) and B(32)) xor (A(14) and B(31)) xor (A(15) and B(30)) xor (A(16) and B(29)) xor (A(17) and B(28)) xor (A(18) and B(27)) xor (A(19) and B(26)) xor (A(20) and B(25)) xor (A(21) and B(24)) xor (A(23) and B(23)) xor (A(23) and B(23)) xor (A(24) and B(21)) xor (A(25) and B(20)) xor (A(26) and B(19)) xor (A(27) and B(18)) xor (A(28) and B(17)) xor (A(29) and B(16)) xor (A(30) and B(15)) xor (A(31) and B(14)) xor (A(32) and B(13)) xor (A(33) and B(12)) xor (A(34) and B(11)) xor (A(35) and B(10)) xor (A(36) and B(9)) xor (A(37) and B(8)) xor (A(38) and B(7)) xor (A(39) and B(6)) xor (A(40) and B(5)) xor (A(41) and B(4)) xor (A(42) and B(3)) xor (A(43) and B(2)) xor (A(44) and B(1)) xor (A(45) and B(0)) xor (A(38) and B(127)) xor (A(39) and B(126)) xor (A(40) and B(125)) xor (A(41) and B(124)) xor (A(42) and B(123)) xor (A(43) and B(122)) xor (A(44) and B(121)) xor (A(45) and B(120)) xor (A(46) and B(119)) xor (A(47) and B(118)) xor (A(48) and B(117)) xor (A(49) and B(116)) xor (A(50) and B(115)) xor (A(51) and B(114)) xor (A(52) and B(113)) xor (A(53) and B(112)) xor (A(54) and B(111)) xor (A(55) and B(110)) xor (A(56) and B(109)) xor (A(57) and B(108)) xor (A(58) and B(107)) xor (A(59) and B(106)) xor (A(60) and B(105)) xor (A(61) and B(104)) xor (A(62) and B(103)) xor (A(63) and B(102)) xor (A(64) and B(101)) xor (A(65) and B(100)) xor (A(66) and B(99)) xor (A(67) and B(98)) xor (A(68) and B(97)) xor (A(69) and B(96)) xor (A(70) and B(95)) xor (A(71) and B(94)) xor (A(72) and B(93)) xor (A(73) and B(92)) xor (A(74) and B(91)) xor (A(75) and B(90)) xor (A(76) and B(89)) xor (A(77) and B(88)) xor (A(78) and B(87)) xor (A(79) and B(86)) xor (A(80) and B(85)) xor (A(81) and B(84)) xor (A(82) and B(83)) xor (A(83) and B(82)) xor (A(84) and B(81)) xor (A(85) and B(80)) xor (A(86) and B(79)) xor (A(87) and B(78)) xor (A(88) and B(77)) xor (A(89) and B(76)) xor (A(90) and B(75)) xor (A(91) and B(74)) xor (A(92) and B(73)) xor (A(93) and B(72)) xor (A(94) and B(71)) xor (A(95) and B(70)) xor (A(96) and B(69)) xor (A(97) and B(68)) xor (A(98) and B(67)) xor (A(99) and B(66)) xor (A(100) and B(65)) xor (A(101) and B(64)) xor (A(102) and B(63)) xor (A(103) and B(62)) xor (A(104) and B(61)) xor (A(105) and B(60)) xor (A(106) and B(59)) xor (A(107) and B(58)) xor (A(108) and B(57)) xor (A(109) and B(56)) xor (A(110) and B(55)) xor (A(111) and B(54)) xor (A(112) and B(53)) xor (A(113) and B(52)) xor (A(114) and B(51)) xor (A(115) and B(50)) xor (A(116) and B(49)) xor (A(117) and B(48)) xor (A(118) and B(47)) xor (A(119) and B(46)) xor (A(120) and B(45)) xor (A(121) and B(44)) xor (A(122) and B(43)) xor (A(123) and B(42)) xor (A(124) and B(41)) xor (A(125) and B(40)) xor (A(126) and B(39)) xor (A(43) and B(127)) xor (A(44) and B(126)) xor (A(45) and B(125)) xor (A(46) and B(124)) xor (A(47) and B(123)) xor (A(48) and B(122)) xor (A(49) and B(121)) xor (A(50) and B(120)) xor (A(51) and B(119)) xor (A(52) and B(118)) xor (A(53) and B(117)) xor (A(54) and B(116)) xor (A(55) and B(115)) xor (A(56) and B(114)) xor (A(57) and B(113)) xor (A(58) and B(112)) xor (A(59) and B(111)) xor (A(60) and B(110)) xor (A(61) and B(109)) xor (A(62) and B(108)) xor (A(63) and B(107)) xor (A(64) and B(106)) xor (A(65) and B(105)) xor (A(66) and B(104)) xor (A(67) and B(103)) xor (A(68) and B(102)) xor (A(69) and B(101)) xor (A(70) and B(100)) xor (A(71) and B(99)) xor (A(72) and B(98)) xor (A(73) and B(97)) xor (A(74) and B(96)) xor (A(75) and B(95)) xor (A(76) and B(94)) xor (A(77) and B(93)) xor (A(78) and B(92)) xor (A(79) and B(91)) xor (A(80) and B(90)) xor (A(81) and B(89)) xor (A(82) and B(88)) xor (A(83) and B(87)) xor (A(84) and B(86)) xor (A(85) and B(85)) xor (A(86) and B(84)) xor (A(87) and B(83)) xor (A(88) and B(82)) xor (A(89) and B(81)) xor (A(90) and B(80)) xor (A(91) and B(79)) xor (A(92) and B(78)) xor (A(93) and B(77)) xor (A(94) and B(76)) xor (A(95) and B(75)) xor (A(96) and B(74)) xor (A(97) and B(73)) xor (A(98) and B(72)) xor (A(99) and B(71)) xor (A(100) and B(70)) xor (A(101) and B(69)) xor (A(102) and B(68)) xor (A(103) and B(67)) xor (A(104) and B(66)) xor (A(105) and B(65)) xor (A(106) and B(64)) xor (A(107) and B(63)) xor (A(108) and B(62)) xor (A(109) and B(61)) xor (A(110) and B(60)) xor (A(111) and B(59)) xor (A(112) and B(58)) xor (A(113) and B(57)) xor (A(114) and B(56)) xor (A(115) and B(55)) xor (A(116) and B(54)) xor (A(117) and B(53)) xor (A(118) and B(52)) xor (A(119) and B(51)) xor (A(120) and B(50)) xor (A(121) and B(49)) xor (A(122) and B(48)) xor (A(123) and B(47)) xor (A(124) and B(46)) xor (A(125) and B(45)) xor (A(126) and B(44)) xor (A(44) and B(127)) xor (A(45) and B(126)) xor (A(46) and B(125)) xor (A(47) and B(124)) xor (A(48) and B(123)) xor (A(49) and B(122)) xor (A(50) and B(121)) xor (A(51) and B(120)) xor (A(52) and B(119)) xor (A(53) and B(118)) xor (A(54) and B(117)) xor (A(55) and B(116)) xor (A(56) and B(115)) xor (A(57) and B(114)) xor (A(58) and B(113)) xor (A(59) and B(112)) xor (A(60) and B(111)) xor (A(61) and B(110)) xor (A(62) and B(109)) xor (A(63) and B(108)) xor (A(64) and B(107)) xor (A(65) and B(106)) xor (A(66) and B(105)) xor (A(67) and B(104)) xor (A(68) and B(103)) xor (A(69) and B(102)) xor (A(70) and B(101)) xor (A(71) and B(100)) xor (A(72) and B(99)) xor (A(73) and B(98)) xor (A(74) and B(97)) xor (A(75) and B(96)) xor (A(76) and B(95)) xor (A(77) and B(94)) xor (A(78) and B(93)) xor (A(79) and B(92)) xor (A(80) and B(91)) xor (A(81) and B(90)) xor (A(82) and B(89)) xor (A(83) and B(88)) xor (A(84) and B(87)) xor (A(85) and B(86)) xor (A(86) and B(85)) xor (A(87) and B(84)) xor (A(88) and B(83)) xor (A(89) and B(82)) xor (A(90) and B(81)) xor (A(91) and B(80)) xor (A(92) and B(79)) xor (A(93) and B(78)) xor (A(94) and B(77)) xor (A(95) and B(76)) xor (A(96) and B(75)) xor (A(97) and B(74)) xor (A(98) and B(73)) xor (A(99) and B(72)) xor (A(100) and B(71)) xor (A(101) and B(70)) xor (A(102) and B(69)) xor (A(103) and B(68)) xor (A(104) and B(67)) xor (A(105) and B(66)) xor (A(106) and B(65)) xor (A(107) and B(64)) xor (A(108) and B(63)) xor (A(109) and B(62)) xor (A(110) and B(61)) xor (A(111) and B(60)) xor (A(112) and B(59)) xor (A(113) and B(58)) xor (A(114) and B(57)) xor (A(115) and B(56)) xor (A(116) and B(55)) xor (A(117) and B(54)) xor (A(118) and B(53)) xor (A(119) and B(52)) xor (A(120) and B(51)) xor (A(121) and B(50)) xor (A(122) and B(49)) xor (A(123) and B(48)) xor (A(124) and B(47)) xor (A(125) and B(46)) xor (A(126) and B(45)) xor (A(45) and B(127)) xor (A(46) and B(126)) xor (A(47) and B(125)) xor (A(48) and B(124)) xor (A(49) and B(123)) xor (A(50) and B(122)) xor (A(51) and B(121)) xor (A(52) and B(120)) xor (A(53) and B(119)) xor (A(54) and B(118)) xor (A(55) and B(117)) xor (A(56) and B(116)) xor (A(57) and B(115)) xor (A(58) and B(114)) xor (A(59) and B(113)) xor (A(60) and B(112)) xor (A(61) and B(111)) xor (A(62) and B(110)) xor (A(63) and B(109)) xor (A(64) and B(108)) xor (A(65) and B(107)) xor (A(66) and B(106)) xor (A(67) and B(105)) xor (A(68) and B(104)) xor (A(69) and B(103)) xor (A(70) and B(102)) xor (A(71) and B(101)) xor (A(72) and B(100)) xor (A(73) and B(99)) xor (A(74) and B(98)) xor (A(75) and B(97)) xor (A(76) and B(96)) xor (A(77) and B(95)) xor (A(78) and B(94)) xor (A(79) and B(93)) xor (A(80) and B(92)) xor (A(81) and B(91)) xor (A(82) and B(90)) xor (A(83) and B(89)) xor (A(84) and B(88)) xor (A(85) and B(87)) xor (A(86) and B(86)) xor (A(87) and B(85)) xor (A(88) and B(84)) xor (A(89) and B(83)) xor (A(90) and B(82)) xor (A(91) and B(81)) xor (A(92) and B(80)) xor (A(93) and B(79)) xor (A(94) and B(78)) xor (A(95) and B(77)) xor (A(96) and B(76)) xor (A(97) and B(75)) xor (A(98) and B(74)) xor (A(99) and B(73)) xor (A(100) and B(72)) xor (A(101) and B(71)) xor (A(102) and B(70)) xor (A(103) and B(69)) xor (A(104) and B(68)) xor (A(105) and B(67)) xor (A(106) and B(66)) xor (A(107) and B(65)) xor (A(108) and B(64)) xor (A(109) and B(63)) xor (A(110) and B(62)) xor (A(111) and B(61)) xor (A(112) and B(60)) xor (A(113) and B(59)) xor (A(114) and B(58)) xor (A(115) and B(57)) xor (A(116) and B(56)) xor (A(117) and B(55)) xor (A(118) and B(54)) xor (A(119) and B(53)) xor (A(120) and B(52)) xor (A(121) and B(51)) xor (A(122) and B(50)) xor (A(123) and B(49)) xor (A(124) and B(48)) xor (A(125) and B(47)) xor (A(126) and B(47));
    C(46)  <= (A(0) and B(46)) xor (A(1) and B(45)) xor (A(2) and B(44)) xor (A(3) and B(43)) xor (A(4) and B(42)) xor (A(5) and B(41)) xor (A(6) and B(40)) xor (A(7) and B(39)) xor (A(8) and B(38)) xor (A(9) and B(37)) xor (A(10) and B(36)) xor (A(11) and B(35)) xor (A(12) and B(34)) xor (A(13) and B(33)) xor (A(14) and B(32)) xor (A(15) and B(31)) xor (A(16) and B(30)) xor (A(17) and B(29)) xor (A(18) and B(28)) xor (A(19) and B(27)) xor (A(20) and B(26)) xor (A(21) and B(25)) xor (A(23) and B(24)) xor (A(23) and B(23)) xor (A(24) and B(23)) xor (A(25) and B(21)) xor (A(26) and B(20)) xor (A(27) and B(19)) xor (A(28) and B(18)) xor (A(29) and B(17)) xor (A(30) and B(16)) xor (A(31) and B(15)) xor (A(32) and B(14)) xor (A(33) and B(13)) xor (A(34) and B(12)) xor (A(35) and B(11)) xor (A(36) and B(10)) xor (A(37) and B(9)) xor (A(38) and B(8)) xor (A(39) and B(7)) xor (A(40) and B(6)) xor (A(41) and B(5)) xor (A(42) and B(4)) xor (A(43) and B(3)) xor (A(44) and B(2)) xor (A(45) and B(1)) xor (A(46) and B(0)) xor (A(39) and B(127)) xor (A(40) and B(126)) xor (A(41) and B(125)) xor (A(42) and B(124)) xor (A(43) and B(123)) xor (A(44) and B(122)) xor (A(45) and B(121)) xor (A(46) and B(120)) xor (A(47) and B(119)) xor (A(48) and B(118)) xor (A(49) and B(117)) xor (A(50) and B(116)) xor (A(51) and B(115)) xor (A(52) and B(114)) xor (A(53) and B(113)) xor (A(54) and B(112)) xor (A(55) and B(111)) xor (A(56) and B(110)) xor (A(57) and B(109)) xor (A(58) and B(108)) xor (A(59) and B(107)) xor (A(60) and B(106)) xor (A(61) and B(105)) xor (A(62) and B(104)) xor (A(63) and B(103)) xor (A(64) and B(102)) xor (A(65) and B(101)) xor (A(66) and B(100)) xor (A(67) and B(99)) xor (A(68) and B(98)) xor (A(69) and B(97)) xor (A(70) and B(96)) xor (A(71) and B(95)) xor (A(72) and B(94)) xor (A(73) and B(93)) xor (A(74) and B(92)) xor (A(75) and B(91)) xor (A(76) and B(90)) xor (A(77) and B(89)) xor (A(78) and B(88)) xor (A(79) and B(87)) xor (A(80) and B(86)) xor (A(81) and B(85)) xor (A(82) and B(84)) xor (A(83) and B(83)) xor (A(84) and B(82)) xor (A(85) and B(81)) xor (A(86) and B(80)) xor (A(87) and B(79)) xor (A(88) and B(78)) xor (A(89) and B(77)) xor (A(90) and B(76)) xor (A(91) and B(75)) xor (A(92) and B(74)) xor (A(93) and B(73)) xor (A(94) and B(72)) xor (A(95) and B(71)) xor (A(96) and B(70)) xor (A(97) and B(69)) xor (A(98) and B(68)) xor (A(99) and B(67)) xor (A(100) and B(66)) xor (A(101) and B(65)) xor (A(102) and B(64)) xor (A(103) and B(63)) xor (A(104) and B(62)) xor (A(105) and B(61)) xor (A(106) and B(60)) xor (A(107) and B(59)) xor (A(108) and B(58)) xor (A(109) and B(57)) xor (A(110) and B(56)) xor (A(111) and B(55)) xor (A(112) and B(54)) xor (A(113) and B(53)) xor (A(114) and B(52)) xor (A(115) and B(51)) xor (A(116) and B(50)) xor (A(117) and B(49)) xor (A(118) and B(48)) xor (A(119) and B(47)) xor (A(120) and B(46)) xor (A(121) and B(45)) xor (A(122) and B(44)) xor (A(123) and B(43)) xor (A(124) and B(42)) xor (A(125) and B(41)) xor (A(126) and B(40)) xor (A(44) and B(127)) xor (A(45) and B(126)) xor (A(46) and B(125)) xor (A(47) and B(124)) xor (A(48) and B(123)) xor (A(49) and B(122)) xor (A(50) and B(121)) xor (A(51) and B(120)) xor (A(52) and B(119)) xor (A(53) and B(118)) xor (A(54) and B(117)) xor (A(55) and B(116)) xor (A(56) and B(115)) xor (A(57) and B(114)) xor (A(58) and B(113)) xor (A(59) and B(112)) xor (A(60) and B(111)) xor (A(61) and B(110)) xor (A(62) and B(109)) xor (A(63) and B(108)) xor (A(64) and B(107)) xor (A(65) and B(106)) xor (A(66) and B(105)) xor (A(67) and B(104)) xor (A(68) and B(103)) xor (A(69) and B(102)) xor (A(70) and B(101)) xor (A(71) and B(100)) xor (A(72) and B(99)) xor (A(73) and B(98)) xor (A(74) and B(97)) xor (A(75) and B(96)) xor (A(76) and B(95)) xor (A(77) and B(94)) xor (A(78) and B(93)) xor (A(79) and B(92)) xor (A(80) and B(91)) xor (A(81) and B(90)) xor (A(82) and B(89)) xor (A(83) and B(88)) xor (A(84) and B(87)) xor (A(85) and B(86)) xor (A(86) and B(85)) xor (A(87) and B(84)) xor (A(88) and B(83)) xor (A(89) and B(82)) xor (A(90) and B(81)) xor (A(91) and B(80)) xor (A(92) and B(79)) xor (A(93) and B(78)) xor (A(94) and B(77)) xor (A(95) and B(76)) xor (A(96) and B(75)) xor (A(97) and B(74)) xor (A(98) and B(73)) xor (A(99) and B(72)) xor (A(100) and B(71)) xor (A(101) and B(70)) xor (A(102) and B(69)) xor (A(103) and B(68)) xor (A(104) and B(67)) xor (A(105) and B(66)) xor (A(106) and B(65)) xor (A(107) and B(64)) xor (A(108) and B(63)) xor (A(109) and B(62)) xor (A(110) and B(61)) xor (A(111) and B(60)) xor (A(112) and B(59)) xor (A(113) and B(58)) xor (A(114) and B(57)) xor (A(115) and B(56)) xor (A(116) and B(55)) xor (A(117) and B(54)) xor (A(118) and B(53)) xor (A(119) and B(52)) xor (A(120) and B(51)) xor (A(121) and B(50)) xor (A(122) and B(49)) xor (A(123) and B(48)) xor (A(124) and B(47)) xor (A(125) and B(46)) xor (A(126) and B(45)) xor (A(45) and B(127)) xor (A(46) and B(126)) xor (A(47) and B(125)) xor (A(48) and B(124)) xor (A(49) and B(123)) xor (A(50) and B(122)) xor (A(51) and B(121)) xor (A(52) and B(120)) xor (A(53) and B(119)) xor (A(54) and B(118)) xor (A(55) and B(117)) xor (A(56) and B(116)) xor (A(57) and B(115)) xor (A(58) and B(114)) xor (A(59) and B(113)) xor (A(60) and B(112)) xor (A(61) and B(111)) xor (A(62) and B(110)) xor (A(63) and B(109)) xor (A(64) and B(108)) xor (A(65) and B(107)) xor (A(66) and B(106)) xor (A(67) and B(105)) xor (A(68) and B(104)) xor (A(69) and B(103)) xor (A(70) and B(102)) xor (A(71) and B(101)) xor (A(72) and B(100)) xor (A(73) and B(99)) xor (A(74) and B(98)) xor (A(75) and B(97)) xor (A(76) and B(96)) xor (A(77) and B(95)) xor (A(78) and B(94)) xor (A(79) and B(93)) xor (A(80) and B(92)) xor (A(81) and B(91)) xor (A(82) and B(90)) xor (A(83) and B(89)) xor (A(84) and B(88)) xor (A(85) and B(87)) xor (A(86) and B(86)) xor (A(87) and B(85)) xor (A(88) and B(84)) xor (A(89) and B(83)) xor (A(90) and B(82)) xor (A(91) and B(81)) xor (A(92) and B(80)) xor (A(93) and B(79)) xor (A(94) and B(78)) xor (A(95) and B(77)) xor (A(96) and B(76)) xor (A(97) and B(75)) xor (A(98) and B(74)) xor (A(99) and B(73)) xor (A(100) and B(72)) xor (A(101) and B(71)) xor (A(102) and B(70)) xor (A(103) and B(69)) xor (A(104) and B(68)) xor (A(105) and B(67)) xor (A(106) and B(66)) xor (A(107) and B(65)) xor (A(108) and B(64)) xor (A(109) and B(63)) xor (A(110) and B(62)) xor (A(111) and B(61)) xor (A(112) and B(60)) xor (A(113) and B(59)) xor (A(114) and B(58)) xor (A(115) and B(57)) xor (A(116) and B(56)) xor (A(117) and B(55)) xor (A(118) and B(54)) xor (A(119) and B(53)) xor (A(120) and B(52)) xor (A(121) and B(51)) xor (A(122) and B(50)) xor (A(123) and B(49)) xor (A(124) and B(48)) xor (A(125) and B(47)) xor (A(126) and B(46)) xor (A(46) and B(127)) xor (A(47) and B(126)) xor (A(48) and B(125)) xor (A(49) and B(124)) xor (A(50) and B(123)) xor (A(51) and B(122)) xor (A(52) and B(121)) xor (A(53) and B(120)) xor (A(54) and B(119)) xor (A(55) and B(118)) xor (A(56) and B(117)) xor (A(57) and B(116)) xor (A(58) and B(115)) xor (A(59) and B(114)) xor (A(60) and B(113)) xor (A(61) and B(112)) xor (A(62) and B(111)) xor (A(63) and B(110)) xor (A(64) and B(109)) xor (A(65) and B(108)) xor (A(66) and B(107)) xor (A(67) and B(106)) xor (A(68) and B(105)) xor (A(69) and B(104)) xor (A(70) and B(103)) xor (A(71) and B(102)) xor (A(72) and B(101)) xor (A(73) and B(100)) xor (A(74) and B(99)) xor (A(75) and B(98)) xor (A(76) and B(97)) xor (A(77) and B(96)) xor (A(78) and B(95)) xor (A(79) and B(94)) xor (A(80) and B(93)) xor (A(81) and B(92)) xor (A(82) and B(91)) xor (A(83) and B(90)) xor (A(84) and B(89)) xor (A(85) and B(88)) xor (A(86) and B(87)) xor (A(87) and B(86)) xor (A(88) and B(85)) xor (A(89) and B(84)) xor (A(90) and B(83)) xor (A(91) and B(82)) xor (A(92) and B(81)) xor (A(93) and B(80)) xor (A(94) and B(79)) xor (A(95) and B(78)) xor (A(96) and B(77)) xor (A(97) and B(76)) xor (A(98) and B(75)) xor (A(99) and B(74)) xor (A(100) and B(73)) xor (A(101) and B(72)) xor (A(102) and B(71)) xor (A(103) and B(70)) xor (A(104) and B(69)) xor (A(105) and B(68)) xor (A(106) and B(67)) xor (A(107) and B(66)) xor (A(108) and B(65)) xor (A(109) and B(64)) xor (A(110) and B(63)) xor (A(111) and B(62)) xor (A(112) and B(61)) xor (A(113) and B(60)) xor (A(114) and B(59)) xor (A(115) and B(58)) xor (A(116) and B(57)) xor (A(117) and B(56)) xor (A(118) and B(55)) xor (A(119) and B(54)) xor (A(120) and B(53)) xor (A(121) and B(52)) xor (A(122) and B(51)) xor (A(123) and B(50)) xor (A(124) and B(49)) xor (A(125) and B(48)) xor (A(126) and B(48));
    C(47)  <= (A(0) and B(47)) xor (A(1) and B(46)) xor (A(2) and B(45)) xor (A(3) and B(44)) xor (A(4) and B(43)) xor (A(5) and B(42)) xor (A(6) and B(41)) xor (A(7) and B(40)) xor (A(8) and B(39)) xor (A(9) and B(38)) xor (A(10) and B(37)) xor (A(11) and B(36)) xor (A(12) and B(35)) xor (A(13) and B(34)) xor (A(14) and B(33)) xor (A(15) and B(32)) xor (A(16) and B(31)) xor (A(17) and B(30)) xor (A(18) and B(29)) xor (A(19) and B(28)) xor (A(20) and B(27)) xor (A(21) and B(26)) xor (A(23) and B(25)) xor (A(23) and B(24)) xor (A(24) and B(23)) xor (A(25) and B(23)) xor (A(26) and B(21)) xor (A(27) and B(20)) xor (A(28) and B(19)) xor (A(29) and B(18)) xor (A(30) and B(17)) xor (A(31) and B(16)) xor (A(32) and B(15)) xor (A(33) and B(14)) xor (A(34) and B(13)) xor (A(35) and B(12)) xor (A(36) and B(11)) xor (A(37) and B(10)) xor (A(38) and B(9)) xor (A(39) and B(8)) xor (A(40) and B(7)) xor (A(41) and B(6)) xor (A(42) and B(5)) xor (A(43) and B(4)) xor (A(44) and B(3)) xor (A(45) and B(2)) xor (A(46) and B(1)) xor (A(47) and B(0)) xor (A(40) and B(127)) xor (A(41) and B(126)) xor (A(42) and B(125)) xor (A(43) and B(124)) xor (A(44) and B(123)) xor (A(45) and B(122)) xor (A(46) and B(121)) xor (A(47) and B(120)) xor (A(48) and B(119)) xor (A(49) and B(118)) xor (A(50) and B(117)) xor (A(51) and B(116)) xor (A(52) and B(115)) xor (A(53) and B(114)) xor (A(54) and B(113)) xor (A(55) and B(112)) xor (A(56) and B(111)) xor (A(57) and B(110)) xor (A(58) and B(109)) xor (A(59) and B(108)) xor (A(60) and B(107)) xor (A(61) and B(106)) xor (A(62) and B(105)) xor (A(63) and B(104)) xor (A(64) and B(103)) xor (A(65) and B(102)) xor (A(66) and B(101)) xor (A(67) and B(100)) xor (A(68) and B(99)) xor (A(69) and B(98)) xor (A(70) and B(97)) xor (A(71) and B(96)) xor (A(72) and B(95)) xor (A(73) and B(94)) xor (A(74) and B(93)) xor (A(75) and B(92)) xor (A(76) and B(91)) xor (A(77) and B(90)) xor (A(78) and B(89)) xor (A(79) and B(88)) xor (A(80) and B(87)) xor (A(81) and B(86)) xor (A(82) and B(85)) xor (A(83) and B(84)) xor (A(84) and B(83)) xor (A(85) and B(82)) xor (A(86) and B(81)) xor (A(87) and B(80)) xor (A(88) and B(79)) xor (A(89) and B(78)) xor (A(90) and B(77)) xor (A(91) and B(76)) xor (A(92) and B(75)) xor (A(93) and B(74)) xor (A(94) and B(73)) xor (A(95) and B(72)) xor (A(96) and B(71)) xor (A(97) and B(70)) xor (A(98) and B(69)) xor (A(99) and B(68)) xor (A(100) and B(67)) xor (A(101) and B(66)) xor (A(102) and B(65)) xor (A(103) and B(64)) xor (A(104) and B(63)) xor (A(105) and B(62)) xor (A(106) and B(61)) xor (A(107) and B(60)) xor (A(108) and B(59)) xor (A(109) and B(58)) xor (A(110) and B(57)) xor (A(111) and B(56)) xor (A(112) and B(55)) xor (A(113) and B(54)) xor (A(114) and B(53)) xor (A(115) and B(52)) xor (A(116) and B(51)) xor (A(117) and B(50)) xor (A(118) and B(49)) xor (A(119) and B(48)) xor (A(120) and B(47)) xor (A(121) and B(46)) xor (A(122) and B(45)) xor (A(123) and B(44)) xor (A(124) and B(43)) xor (A(125) and B(42)) xor (A(126) and B(41)) xor (A(45) and B(127)) xor (A(46) and B(126)) xor (A(47) and B(125)) xor (A(48) and B(124)) xor (A(49) and B(123)) xor (A(50) and B(122)) xor (A(51) and B(121)) xor (A(52) and B(120)) xor (A(53) and B(119)) xor (A(54) and B(118)) xor (A(55) and B(117)) xor (A(56) and B(116)) xor (A(57) and B(115)) xor (A(58) and B(114)) xor (A(59) and B(113)) xor (A(60) and B(112)) xor (A(61) and B(111)) xor (A(62) and B(110)) xor (A(63) and B(109)) xor (A(64) and B(108)) xor (A(65) and B(107)) xor (A(66) and B(106)) xor (A(67) and B(105)) xor (A(68) and B(104)) xor (A(69) and B(103)) xor (A(70) and B(102)) xor (A(71) and B(101)) xor (A(72) and B(100)) xor (A(73) and B(99)) xor (A(74) and B(98)) xor (A(75) and B(97)) xor (A(76) and B(96)) xor (A(77) and B(95)) xor (A(78) and B(94)) xor (A(79) and B(93)) xor (A(80) and B(92)) xor (A(81) and B(91)) xor (A(82) and B(90)) xor (A(83) and B(89)) xor (A(84) and B(88)) xor (A(85) and B(87)) xor (A(86) and B(86)) xor (A(87) and B(85)) xor (A(88) and B(84)) xor (A(89) and B(83)) xor (A(90) and B(82)) xor (A(91) and B(81)) xor (A(92) and B(80)) xor (A(93) and B(79)) xor (A(94) and B(78)) xor (A(95) and B(77)) xor (A(96) and B(76)) xor (A(97) and B(75)) xor (A(98) and B(74)) xor (A(99) and B(73)) xor (A(100) and B(72)) xor (A(101) and B(71)) xor (A(102) and B(70)) xor (A(103) and B(69)) xor (A(104) and B(68)) xor (A(105) and B(67)) xor (A(106) and B(66)) xor (A(107) and B(65)) xor (A(108) and B(64)) xor (A(109) and B(63)) xor (A(110) and B(62)) xor (A(111) and B(61)) xor (A(112) and B(60)) xor (A(113) and B(59)) xor (A(114) and B(58)) xor (A(115) and B(57)) xor (A(116) and B(56)) xor (A(117) and B(55)) xor (A(118) and B(54)) xor (A(119) and B(53)) xor (A(120) and B(52)) xor (A(121) and B(51)) xor (A(122) and B(50)) xor (A(123) and B(49)) xor (A(124) and B(48)) xor (A(125) and B(47)) xor (A(126) and B(46)) xor (A(46) and B(127)) xor (A(47) and B(126)) xor (A(48) and B(125)) xor (A(49) and B(124)) xor (A(50) and B(123)) xor (A(51) and B(122)) xor (A(52) and B(121)) xor (A(53) and B(120)) xor (A(54) and B(119)) xor (A(55) and B(118)) xor (A(56) and B(117)) xor (A(57) and B(116)) xor (A(58) and B(115)) xor (A(59) and B(114)) xor (A(60) and B(113)) xor (A(61) and B(112)) xor (A(62) and B(111)) xor (A(63) and B(110)) xor (A(64) and B(109)) xor (A(65) and B(108)) xor (A(66) and B(107)) xor (A(67) and B(106)) xor (A(68) and B(105)) xor (A(69) and B(104)) xor (A(70) and B(103)) xor (A(71) and B(102)) xor (A(72) and B(101)) xor (A(73) and B(100)) xor (A(74) and B(99)) xor (A(75) and B(98)) xor (A(76) and B(97)) xor (A(77) and B(96)) xor (A(78) and B(95)) xor (A(79) and B(94)) xor (A(80) and B(93)) xor (A(81) and B(92)) xor (A(82) and B(91)) xor (A(83) and B(90)) xor (A(84) and B(89)) xor (A(85) and B(88)) xor (A(86) and B(87)) xor (A(87) and B(86)) xor (A(88) and B(85)) xor (A(89) and B(84)) xor (A(90) and B(83)) xor (A(91) and B(82)) xor (A(92) and B(81)) xor (A(93) and B(80)) xor (A(94) and B(79)) xor (A(95) and B(78)) xor (A(96) and B(77)) xor (A(97) and B(76)) xor (A(98) and B(75)) xor (A(99) and B(74)) xor (A(100) and B(73)) xor (A(101) and B(72)) xor (A(102) and B(71)) xor (A(103) and B(70)) xor (A(104) and B(69)) xor (A(105) and B(68)) xor (A(106) and B(67)) xor (A(107) and B(66)) xor (A(108) and B(65)) xor (A(109) and B(64)) xor (A(110) and B(63)) xor (A(111) and B(62)) xor (A(112) and B(61)) xor (A(113) and B(60)) xor (A(114) and B(59)) xor (A(115) and B(58)) xor (A(116) and B(57)) xor (A(117) and B(56)) xor (A(118) and B(55)) xor (A(119) and B(54)) xor (A(120) and B(53)) xor (A(121) and B(52)) xor (A(122) and B(51)) xor (A(123) and B(50)) xor (A(124) and B(49)) xor (A(125) and B(48)) xor (A(126) and B(47)) xor (A(47) and B(127)) xor (A(48) and B(126)) xor (A(49) and B(125)) xor (A(50) and B(124)) xor (A(51) and B(123)) xor (A(52) and B(122)) xor (A(53) and B(121)) xor (A(54) and B(120)) xor (A(55) and B(119)) xor (A(56) and B(118)) xor (A(57) and B(117)) xor (A(58) and B(116)) xor (A(59) and B(115)) xor (A(60) and B(114)) xor (A(61) and B(113)) xor (A(62) and B(112)) xor (A(63) and B(111)) xor (A(64) and B(110)) xor (A(65) and B(109)) xor (A(66) and B(108)) xor (A(67) and B(107)) xor (A(68) and B(106)) xor (A(69) and B(105)) xor (A(70) and B(104)) xor (A(71) and B(103)) xor (A(72) and B(102)) xor (A(73) and B(101)) xor (A(74) and B(100)) xor (A(75) and B(99)) xor (A(76) and B(98)) xor (A(77) and B(97)) xor (A(78) and B(96)) xor (A(79) and B(95)) xor (A(80) and B(94)) xor (A(81) and B(93)) xor (A(82) and B(92)) xor (A(83) and B(91)) xor (A(84) and B(90)) xor (A(85) and B(89)) xor (A(86) and B(88)) xor (A(87) and B(87)) xor (A(88) and B(86)) xor (A(89) and B(85)) xor (A(90) and B(84)) xor (A(91) and B(83)) xor (A(92) and B(82)) xor (A(93) and B(81)) xor (A(94) and B(80)) xor (A(95) and B(79)) xor (A(96) and B(78)) xor (A(97) and B(77)) xor (A(98) and B(76)) xor (A(99) and B(75)) xor (A(100) and B(74)) xor (A(101) and B(73)) xor (A(102) and B(72)) xor (A(103) and B(71)) xor (A(104) and B(70)) xor (A(105) and B(69)) xor (A(106) and B(68)) xor (A(107) and B(67)) xor (A(108) and B(66)) xor (A(109) and B(65)) xor (A(110) and B(64)) xor (A(111) and B(63)) xor (A(112) and B(62)) xor (A(113) and B(61)) xor (A(114) and B(60)) xor (A(115) and B(59)) xor (A(116) and B(58)) xor (A(117) and B(57)) xor (A(118) and B(56)) xor (A(119) and B(55)) xor (A(120) and B(54)) xor (A(121) and B(53)) xor (A(122) and B(52)) xor (A(123) and B(51)) xor (A(124) and B(50)) xor (A(125) and B(49)) xor (A(126) and B(49));
    C(48)  <= (A(0) and B(48)) xor (A(1) and B(47)) xor (A(2) and B(46)) xor (A(3) and B(45)) xor (A(4) and B(44)) xor (A(5) and B(43)) xor (A(6) and B(42)) xor (A(7) and B(41)) xor (A(8) and B(40)) xor (A(9) and B(39)) xor (A(10) and B(38)) xor (A(11) and B(37)) xor (A(12) and B(36)) xor (A(13) and B(35)) xor (A(14) and B(34)) xor (A(15) and B(33)) xor (A(16) and B(32)) xor (A(17) and B(31)) xor (A(18) and B(30)) xor (A(19) and B(29)) xor (A(20) and B(28)) xor (A(21) and B(27)) xor (A(23) and B(26)) xor (A(23) and B(25)) xor (A(24) and B(24)) xor (A(25) and B(23)) xor (A(26) and B(23)) xor (A(27) and B(21)) xor (A(28) and B(20)) xor (A(29) and B(19)) xor (A(30) and B(18)) xor (A(31) and B(17)) xor (A(32) and B(16)) xor (A(33) and B(15)) xor (A(34) and B(14)) xor (A(35) and B(13)) xor (A(36) and B(12)) xor (A(37) and B(11)) xor (A(38) and B(10)) xor (A(39) and B(9)) xor (A(40) and B(8)) xor (A(41) and B(7)) xor (A(42) and B(6)) xor (A(43) and B(5)) xor (A(44) and B(4)) xor (A(45) and B(3)) xor (A(46) and B(2)) xor (A(47) and B(1)) xor (A(48) and B(0)) xor (A(41) and B(127)) xor (A(42) and B(126)) xor (A(43) and B(125)) xor (A(44) and B(124)) xor (A(45) and B(123)) xor (A(46) and B(122)) xor (A(47) and B(121)) xor (A(48) and B(120)) xor (A(49) and B(119)) xor (A(50) and B(118)) xor (A(51) and B(117)) xor (A(52) and B(116)) xor (A(53) and B(115)) xor (A(54) and B(114)) xor (A(55) and B(113)) xor (A(56) and B(112)) xor (A(57) and B(111)) xor (A(58) and B(110)) xor (A(59) and B(109)) xor (A(60) and B(108)) xor (A(61) and B(107)) xor (A(62) and B(106)) xor (A(63) and B(105)) xor (A(64) and B(104)) xor (A(65) and B(103)) xor (A(66) and B(102)) xor (A(67) and B(101)) xor (A(68) and B(100)) xor (A(69) and B(99)) xor (A(70) and B(98)) xor (A(71) and B(97)) xor (A(72) and B(96)) xor (A(73) and B(95)) xor (A(74) and B(94)) xor (A(75) and B(93)) xor (A(76) and B(92)) xor (A(77) and B(91)) xor (A(78) and B(90)) xor (A(79) and B(89)) xor (A(80) and B(88)) xor (A(81) and B(87)) xor (A(82) and B(86)) xor (A(83) and B(85)) xor (A(84) and B(84)) xor (A(85) and B(83)) xor (A(86) and B(82)) xor (A(87) and B(81)) xor (A(88) and B(80)) xor (A(89) and B(79)) xor (A(90) and B(78)) xor (A(91) and B(77)) xor (A(92) and B(76)) xor (A(93) and B(75)) xor (A(94) and B(74)) xor (A(95) and B(73)) xor (A(96) and B(72)) xor (A(97) and B(71)) xor (A(98) and B(70)) xor (A(99) and B(69)) xor (A(100) and B(68)) xor (A(101) and B(67)) xor (A(102) and B(66)) xor (A(103) and B(65)) xor (A(104) and B(64)) xor (A(105) and B(63)) xor (A(106) and B(62)) xor (A(107) and B(61)) xor (A(108) and B(60)) xor (A(109) and B(59)) xor (A(110) and B(58)) xor (A(111) and B(57)) xor (A(112) and B(56)) xor (A(113) and B(55)) xor (A(114) and B(54)) xor (A(115) and B(53)) xor (A(116) and B(52)) xor (A(117) and B(51)) xor (A(118) and B(50)) xor (A(119) and B(49)) xor (A(120) and B(48)) xor (A(121) and B(47)) xor (A(122) and B(46)) xor (A(123) and B(45)) xor (A(124) and B(44)) xor (A(125) and B(43)) xor (A(126) and B(42)) xor (A(46) and B(127)) xor (A(47) and B(126)) xor (A(48) and B(125)) xor (A(49) and B(124)) xor (A(50) and B(123)) xor (A(51) and B(122)) xor (A(52) and B(121)) xor (A(53) and B(120)) xor (A(54) and B(119)) xor (A(55) and B(118)) xor (A(56) and B(117)) xor (A(57) and B(116)) xor (A(58) and B(115)) xor (A(59) and B(114)) xor (A(60) and B(113)) xor (A(61) and B(112)) xor (A(62) and B(111)) xor (A(63) and B(110)) xor (A(64) and B(109)) xor (A(65) and B(108)) xor (A(66) and B(107)) xor (A(67) and B(106)) xor (A(68) and B(105)) xor (A(69) and B(104)) xor (A(70) and B(103)) xor (A(71) and B(102)) xor (A(72) and B(101)) xor (A(73) and B(100)) xor (A(74) and B(99)) xor (A(75) and B(98)) xor (A(76) and B(97)) xor (A(77) and B(96)) xor (A(78) and B(95)) xor (A(79) and B(94)) xor (A(80) and B(93)) xor (A(81) and B(92)) xor (A(82) and B(91)) xor (A(83) and B(90)) xor (A(84) and B(89)) xor (A(85) and B(88)) xor (A(86) and B(87)) xor (A(87) and B(86)) xor (A(88) and B(85)) xor (A(89) and B(84)) xor (A(90) and B(83)) xor (A(91) and B(82)) xor (A(92) and B(81)) xor (A(93) and B(80)) xor (A(94) and B(79)) xor (A(95) and B(78)) xor (A(96) and B(77)) xor (A(97) and B(76)) xor (A(98) and B(75)) xor (A(99) and B(74)) xor (A(100) and B(73)) xor (A(101) and B(72)) xor (A(102) and B(71)) xor (A(103) and B(70)) xor (A(104) and B(69)) xor (A(105) and B(68)) xor (A(106) and B(67)) xor (A(107) and B(66)) xor (A(108) and B(65)) xor (A(109) and B(64)) xor (A(110) and B(63)) xor (A(111) and B(62)) xor (A(112) and B(61)) xor (A(113) and B(60)) xor (A(114) and B(59)) xor (A(115) and B(58)) xor (A(116) and B(57)) xor (A(117) and B(56)) xor (A(118) and B(55)) xor (A(119) and B(54)) xor (A(120) and B(53)) xor (A(121) and B(52)) xor (A(122) and B(51)) xor (A(123) and B(50)) xor (A(124) and B(49)) xor (A(125) and B(48)) xor (A(126) and B(47)) xor (A(47) and B(127)) xor (A(48) and B(126)) xor (A(49) and B(125)) xor (A(50) and B(124)) xor (A(51) and B(123)) xor (A(52) and B(122)) xor (A(53) and B(121)) xor (A(54) and B(120)) xor (A(55) and B(119)) xor (A(56) and B(118)) xor (A(57) and B(117)) xor (A(58) and B(116)) xor (A(59) and B(115)) xor (A(60) and B(114)) xor (A(61) and B(113)) xor (A(62) and B(112)) xor (A(63) and B(111)) xor (A(64) and B(110)) xor (A(65) and B(109)) xor (A(66) and B(108)) xor (A(67) and B(107)) xor (A(68) and B(106)) xor (A(69) and B(105)) xor (A(70) and B(104)) xor (A(71) and B(103)) xor (A(72) and B(102)) xor (A(73) and B(101)) xor (A(74) and B(100)) xor (A(75) and B(99)) xor (A(76) and B(98)) xor (A(77) and B(97)) xor (A(78) and B(96)) xor (A(79) and B(95)) xor (A(80) and B(94)) xor (A(81) and B(93)) xor (A(82) and B(92)) xor (A(83) and B(91)) xor (A(84) and B(90)) xor (A(85) and B(89)) xor (A(86) and B(88)) xor (A(87) and B(87)) xor (A(88) and B(86)) xor (A(89) and B(85)) xor (A(90) and B(84)) xor (A(91) and B(83)) xor (A(92) and B(82)) xor (A(93) and B(81)) xor (A(94) and B(80)) xor (A(95) and B(79)) xor (A(96) and B(78)) xor (A(97) and B(77)) xor (A(98) and B(76)) xor (A(99) and B(75)) xor (A(100) and B(74)) xor (A(101) and B(73)) xor (A(102) and B(72)) xor (A(103) and B(71)) xor (A(104) and B(70)) xor (A(105) and B(69)) xor (A(106) and B(68)) xor (A(107) and B(67)) xor (A(108) and B(66)) xor (A(109) and B(65)) xor (A(110) and B(64)) xor (A(111) and B(63)) xor (A(112) and B(62)) xor (A(113) and B(61)) xor (A(114) and B(60)) xor (A(115) and B(59)) xor (A(116) and B(58)) xor (A(117) and B(57)) xor (A(118) and B(56)) xor (A(119) and B(55)) xor (A(120) and B(54)) xor (A(121) and B(53)) xor (A(122) and B(52)) xor (A(123) and B(51)) xor (A(124) and B(50)) xor (A(125) and B(49)) xor (A(126) and B(48)) xor (A(48) and B(127)) xor (A(49) and B(126)) xor (A(50) and B(125)) xor (A(51) and B(124)) xor (A(52) and B(123)) xor (A(53) and B(122)) xor (A(54) and B(121)) xor (A(55) and B(120)) xor (A(56) and B(119)) xor (A(57) and B(118)) xor (A(58) and B(117)) xor (A(59) and B(116)) xor (A(60) and B(115)) xor (A(61) and B(114)) xor (A(62) and B(113)) xor (A(63) and B(112)) xor (A(64) and B(111)) xor (A(65) and B(110)) xor (A(66) and B(109)) xor (A(67) and B(108)) xor (A(68) and B(107)) xor (A(69) and B(106)) xor (A(70) and B(105)) xor (A(71) and B(104)) xor (A(72) and B(103)) xor (A(73) and B(102)) xor (A(74) and B(101)) xor (A(75) and B(100)) xor (A(76) and B(99)) xor (A(77) and B(98)) xor (A(78) and B(97)) xor (A(79) and B(96)) xor (A(80) and B(95)) xor (A(81) and B(94)) xor (A(82) and B(93)) xor (A(83) and B(92)) xor (A(84) and B(91)) xor (A(85) and B(90)) xor (A(86) and B(89)) xor (A(87) and B(88)) xor (A(88) and B(87)) xor (A(89) and B(86)) xor (A(90) and B(85)) xor (A(91) and B(84)) xor (A(92) and B(83)) xor (A(93) and B(82)) xor (A(94) and B(81)) xor (A(95) and B(80)) xor (A(96) and B(79)) xor (A(97) and B(78)) xor (A(98) and B(77)) xor (A(99) and B(76)) xor (A(100) and B(75)) xor (A(101) and B(74)) xor (A(102) and B(73)) xor (A(103) and B(72)) xor (A(104) and B(71)) xor (A(105) and B(70)) xor (A(106) and B(69)) xor (A(107) and B(68)) xor (A(108) and B(67)) xor (A(109) and B(66)) xor (A(110) and B(65)) xor (A(111) and B(64)) xor (A(112) and B(63)) xor (A(113) and B(62)) xor (A(114) and B(61)) xor (A(115) and B(60)) xor (A(116) and B(59)) xor (A(117) and B(58)) xor (A(118) and B(57)) xor (A(119) and B(56)) xor (A(120) and B(55)) xor (A(121) and B(54)) xor (A(122) and B(53)) xor (A(123) and B(52)) xor (A(124) and B(51)) xor (A(125) and B(50)) xor (A(126) and B(50));
    C(49)  <= (A(0) and B(49)) xor (A(1) and B(48)) xor (A(2) and B(47)) xor (A(3) and B(46)) xor (A(4) and B(45)) xor (A(5) and B(44)) xor (A(6) and B(43)) xor (A(7) and B(42)) xor (A(8) and B(41)) xor (A(9) and B(40)) xor (A(10) and B(39)) xor (A(11) and B(38)) xor (A(12) and B(37)) xor (A(13) and B(36)) xor (A(14) and B(35)) xor (A(15) and B(34)) xor (A(16) and B(33)) xor (A(17) and B(32)) xor (A(18) and B(31)) xor (A(19) and B(30)) xor (A(20) and B(29)) xor (A(21) and B(28)) xor (A(23) and B(27)) xor (A(23) and B(26)) xor (A(24) and B(25)) xor (A(25) and B(24)) xor (A(26) and B(23)) xor (A(27) and B(23)) xor (A(28) and B(21)) xor (A(29) and B(20)) xor (A(30) and B(19)) xor (A(31) and B(18)) xor (A(32) and B(17)) xor (A(33) and B(16)) xor (A(34) and B(15)) xor (A(35) and B(14)) xor (A(36) and B(13)) xor (A(37) and B(12)) xor (A(38) and B(11)) xor (A(39) and B(10)) xor (A(40) and B(9)) xor (A(41) and B(8)) xor (A(42) and B(7)) xor (A(43) and B(6)) xor (A(44) and B(5)) xor (A(45) and B(4)) xor (A(46) and B(3)) xor (A(47) and B(2)) xor (A(48) and B(1)) xor (A(49) and B(0)) xor (A(42) and B(127)) xor (A(43) and B(126)) xor (A(44) and B(125)) xor (A(45) and B(124)) xor (A(46) and B(123)) xor (A(47) and B(122)) xor (A(48) and B(121)) xor (A(49) and B(120)) xor (A(50) and B(119)) xor (A(51) and B(118)) xor (A(52) and B(117)) xor (A(53) and B(116)) xor (A(54) and B(115)) xor (A(55) and B(114)) xor (A(56) and B(113)) xor (A(57) and B(112)) xor (A(58) and B(111)) xor (A(59) and B(110)) xor (A(60) and B(109)) xor (A(61) and B(108)) xor (A(62) and B(107)) xor (A(63) and B(106)) xor (A(64) and B(105)) xor (A(65) and B(104)) xor (A(66) and B(103)) xor (A(67) and B(102)) xor (A(68) and B(101)) xor (A(69) and B(100)) xor (A(70) and B(99)) xor (A(71) and B(98)) xor (A(72) and B(97)) xor (A(73) and B(96)) xor (A(74) and B(95)) xor (A(75) and B(94)) xor (A(76) and B(93)) xor (A(77) and B(92)) xor (A(78) and B(91)) xor (A(79) and B(90)) xor (A(80) and B(89)) xor (A(81) and B(88)) xor (A(82) and B(87)) xor (A(83) and B(86)) xor (A(84) and B(85)) xor (A(85) and B(84)) xor (A(86) and B(83)) xor (A(87) and B(82)) xor (A(88) and B(81)) xor (A(89) and B(80)) xor (A(90) and B(79)) xor (A(91) and B(78)) xor (A(92) and B(77)) xor (A(93) and B(76)) xor (A(94) and B(75)) xor (A(95) and B(74)) xor (A(96) and B(73)) xor (A(97) and B(72)) xor (A(98) and B(71)) xor (A(99) and B(70)) xor (A(100) and B(69)) xor (A(101) and B(68)) xor (A(102) and B(67)) xor (A(103) and B(66)) xor (A(104) and B(65)) xor (A(105) and B(64)) xor (A(106) and B(63)) xor (A(107) and B(62)) xor (A(108) and B(61)) xor (A(109) and B(60)) xor (A(110) and B(59)) xor (A(111) and B(58)) xor (A(112) and B(57)) xor (A(113) and B(56)) xor (A(114) and B(55)) xor (A(115) and B(54)) xor (A(116) and B(53)) xor (A(117) and B(52)) xor (A(118) and B(51)) xor (A(119) and B(50)) xor (A(120) and B(49)) xor (A(121) and B(48)) xor (A(122) and B(47)) xor (A(123) and B(46)) xor (A(124) and B(45)) xor (A(125) and B(44)) xor (A(126) and B(43)) xor (A(47) and B(127)) xor (A(48) and B(126)) xor (A(49) and B(125)) xor (A(50) and B(124)) xor (A(51) and B(123)) xor (A(52) and B(122)) xor (A(53) and B(121)) xor (A(54) and B(120)) xor (A(55) and B(119)) xor (A(56) and B(118)) xor (A(57) and B(117)) xor (A(58) and B(116)) xor (A(59) and B(115)) xor (A(60) and B(114)) xor (A(61) and B(113)) xor (A(62) and B(112)) xor (A(63) and B(111)) xor (A(64) and B(110)) xor (A(65) and B(109)) xor (A(66) and B(108)) xor (A(67) and B(107)) xor (A(68) and B(106)) xor (A(69) and B(105)) xor (A(70) and B(104)) xor (A(71) and B(103)) xor (A(72) and B(102)) xor (A(73) and B(101)) xor (A(74) and B(100)) xor (A(75) and B(99)) xor (A(76) and B(98)) xor (A(77) and B(97)) xor (A(78) and B(96)) xor (A(79) and B(95)) xor (A(80) and B(94)) xor (A(81) and B(93)) xor (A(82) and B(92)) xor (A(83) and B(91)) xor (A(84) and B(90)) xor (A(85) and B(89)) xor (A(86) and B(88)) xor (A(87) and B(87)) xor (A(88) and B(86)) xor (A(89) and B(85)) xor (A(90) and B(84)) xor (A(91) and B(83)) xor (A(92) and B(82)) xor (A(93) and B(81)) xor (A(94) and B(80)) xor (A(95) and B(79)) xor (A(96) and B(78)) xor (A(97) and B(77)) xor (A(98) and B(76)) xor (A(99) and B(75)) xor (A(100) and B(74)) xor (A(101) and B(73)) xor (A(102) and B(72)) xor (A(103) and B(71)) xor (A(104) and B(70)) xor (A(105) and B(69)) xor (A(106) and B(68)) xor (A(107) and B(67)) xor (A(108) and B(66)) xor (A(109) and B(65)) xor (A(110) and B(64)) xor (A(111) and B(63)) xor (A(112) and B(62)) xor (A(113) and B(61)) xor (A(114) and B(60)) xor (A(115) and B(59)) xor (A(116) and B(58)) xor (A(117) and B(57)) xor (A(118) and B(56)) xor (A(119) and B(55)) xor (A(120) and B(54)) xor (A(121) and B(53)) xor (A(122) and B(52)) xor (A(123) and B(51)) xor (A(124) and B(50)) xor (A(125) and B(49)) xor (A(126) and B(48)) xor (A(48) and B(127)) xor (A(49) and B(126)) xor (A(50) and B(125)) xor (A(51) and B(124)) xor (A(52) and B(123)) xor (A(53) and B(122)) xor (A(54) and B(121)) xor (A(55) and B(120)) xor (A(56) and B(119)) xor (A(57) and B(118)) xor (A(58) and B(117)) xor (A(59) and B(116)) xor (A(60) and B(115)) xor (A(61) and B(114)) xor (A(62) and B(113)) xor (A(63) and B(112)) xor (A(64) and B(111)) xor (A(65) and B(110)) xor (A(66) and B(109)) xor (A(67) and B(108)) xor (A(68) and B(107)) xor (A(69) and B(106)) xor (A(70) and B(105)) xor (A(71) and B(104)) xor (A(72) and B(103)) xor (A(73) and B(102)) xor (A(74) and B(101)) xor (A(75) and B(100)) xor (A(76) and B(99)) xor (A(77) and B(98)) xor (A(78) and B(97)) xor (A(79) and B(96)) xor (A(80) and B(95)) xor (A(81) and B(94)) xor (A(82) and B(93)) xor (A(83) and B(92)) xor (A(84) and B(91)) xor (A(85) and B(90)) xor (A(86) and B(89)) xor (A(87) and B(88)) xor (A(88) and B(87)) xor (A(89) and B(86)) xor (A(90) and B(85)) xor (A(91) and B(84)) xor (A(92) and B(83)) xor (A(93) and B(82)) xor (A(94) and B(81)) xor (A(95) and B(80)) xor (A(96) and B(79)) xor (A(97) and B(78)) xor (A(98) and B(77)) xor (A(99) and B(76)) xor (A(100) and B(75)) xor (A(101) and B(74)) xor (A(102) and B(73)) xor (A(103) and B(72)) xor (A(104) and B(71)) xor (A(105) and B(70)) xor (A(106) and B(69)) xor (A(107) and B(68)) xor (A(108) and B(67)) xor (A(109) and B(66)) xor (A(110) and B(65)) xor (A(111) and B(64)) xor (A(112) and B(63)) xor (A(113) and B(62)) xor (A(114) and B(61)) xor (A(115) and B(60)) xor (A(116) and B(59)) xor (A(117) and B(58)) xor (A(118) and B(57)) xor (A(119) and B(56)) xor (A(120) and B(55)) xor (A(121) and B(54)) xor (A(122) and B(53)) xor (A(123) and B(52)) xor (A(124) and B(51)) xor (A(125) and B(50)) xor (A(126) and B(49)) xor (A(49) and B(127)) xor (A(50) and B(126)) xor (A(51) and B(125)) xor (A(52) and B(124)) xor (A(53) and B(123)) xor (A(54) and B(122)) xor (A(55) and B(121)) xor (A(56) and B(120)) xor (A(57) and B(119)) xor (A(58) and B(118)) xor (A(59) and B(117)) xor (A(60) and B(116)) xor (A(61) and B(115)) xor (A(62) and B(114)) xor (A(63) and B(113)) xor (A(64) and B(112)) xor (A(65) and B(111)) xor (A(66) and B(110)) xor (A(67) and B(109)) xor (A(68) and B(108)) xor (A(69) and B(107)) xor (A(70) and B(106)) xor (A(71) and B(105)) xor (A(72) and B(104)) xor (A(73) and B(103)) xor (A(74) and B(102)) xor (A(75) and B(101)) xor (A(76) and B(100)) xor (A(77) and B(99)) xor (A(78) and B(98)) xor (A(79) and B(97)) xor (A(80) and B(96)) xor (A(81) and B(95)) xor (A(82) and B(94)) xor (A(83) and B(93)) xor (A(84) and B(92)) xor (A(85) and B(91)) xor (A(86) and B(90)) xor (A(87) and B(89)) xor (A(88) and B(88)) xor (A(89) and B(87)) xor (A(90) and B(86)) xor (A(91) and B(85)) xor (A(92) and B(84)) xor (A(93) and B(83)) xor (A(94) and B(82)) xor (A(95) and B(81)) xor (A(96) and B(80)) xor (A(97) and B(79)) xor (A(98) and B(78)) xor (A(99) and B(77)) xor (A(100) and B(76)) xor (A(101) and B(75)) xor (A(102) and B(74)) xor (A(103) and B(73)) xor (A(104) and B(72)) xor (A(105) and B(71)) xor (A(106) and B(70)) xor (A(107) and B(69)) xor (A(108) and B(68)) xor (A(109) and B(67)) xor (A(110) and B(66)) xor (A(111) and B(65)) xor (A(112) and B(64)) xor (A(113) and B(63)) xor (A(114) and B(62)) xor (A(115) and B(61)) xor (A(116) and B(60)) xor (A(117) and B(59)) xor (A(118) and B(58)) xor (A(119) and B(57)) xor (A(120) and B(56)) xor (A(121) and B(55)) xor (A(122) and B(54)) xor (A(123) and B(53)) xor (A(124) and B(52)) xor (A(125) and B(51)) xor (A(126) and B(51));
    C(50)  <= (A(0) and B(50)) xor (A(1) and B(49)) xor (A(2) and B(48)) xor (A(3) and B(47)) xor (A(4) and B(46)) xor (A(5) and B(45)) xor (A(6) and B(44)) xor (A(7) and B(43)) xor (A(8) and B(42)) xor (A(9) and B(41)) xor (A(10) and B(40)) xor (A(11) and B(39)) xor (A(12) and B(38)) xor (A(13) and B(37)) xor (A(14) and B(36)) xor (A(15) and B(35)) xor (A(16) and B(34)) xor (A(17) and B(33)) xor (A(18) and B(32)) xor (A(19) and B(31)) xor (A(20) and B(30)) xor (A(21) and B(29)) xor (A(23) and B(28)) xor (A(23) and B(27)) xor (A(24) and B(26)) xor (A(25) and B(25)) xor (A(26) and B(24)) xor (A(27) and B(23)) xor (A(28) and B(23)) xor (A(29) and B(21)) xor (A(30) and B(20)) xor (A(31) and B(19)) xor (A(32) and B(18)) xor (A(33) and B(17)) xor (A(34) and B(16)) xor (A(35) and B(15)) xor (A(36) and B(14)) xor (A(37) and B(13)) xor (A(38) and B(12)) xor (A(39) and B(11)) xor (A(40) and B(10)) xor (A(41) and B(9)) xor (A(42) and B(8)) xor (A(43) and B(7)) xor (A(44) and B(6)) xor (A(45) and B(5)) xor (A(46) and B(4)) xor (A(47) and B(3)) xor (A(48) and B(2)) xor (A(49) and B(1)) xor (A(50) and B(0)) xor (A(43) and B(127)) xor (A(44) and B(126)) xor (A(45) and B(125)) xor (A(46) and B(124)) xor (A(47) and B(123)) xor (A(48) and B(122)) xor (A(49) and B(121)) xor (A(50) and B(120)) xor (A(51) and B(119)) xor (A(52) and B(118)) xor (A(53) and B(117)) xor (A(54) and B(116)) xor (A(55) and B(115)) xor (A(56) and B(114)) xor (A(57) and B(113)) xor (A(58) and B(112)) xor (A(59) and B(111)) xor (A(60) and B(110)) xor (A(61) and B(109)) xor (A(62) and B(108)) xor (A(63) and B(107)) xor (A(64) and B(106)) xor (A(65) and B(105)) xor (A(66) and B(104)) xor (A(67) and B(103)) xor (A(68) and B(102)) xor (A(69) and B(101)) xor (A(70) and B(100)) xor (A(71) and B(99)) xor (A(72) and B(98)) xor (A(73) and B(97)) xor (A(74) and B(96)) xor (A(75) and B(95)) xor (A(76) and B(94)) xor (A(77) and B(93)) xor (A(78) and B(92)) xor (A(79) and B(91)) xor (A(80) and B(90)) xor (A(81) and B(89)) xor (A(82) and B(88)) xor (A(83) and B(87)) xor (A(84) and B(86)) xor (A(85) and B(85)) xor (A(86) and B(84)) xor (A(87) and B(83)) xor (A(88) and B(82)) xor (A(89) and B(81)) xor (A(90) and B(80)) xor (A(91) and B(79)) xor (A(92) and B(78)) xor (A(93) and B(77)) xor (A(94) and B(76)) xor (A(95) and B(75)) xor (A(96) and B(74)) xor (A(97) and B(73)) xor (A(98) and B(72)) xor (A(99) and B(71)) xor (A(100) and B(70)) xor (A(101) and B(69)) xor (A(102) and B(68)) xor (A(103) and B(67)) xor (A(104) and B(66)) xor (A(105) and B(65)) xor (A(106) and B(64)) xor (A(107) and B(63)) xor (A(108) and B(62)) xor (A(109) and B(61)) xor (A(110) and B(60)) xor (A(111) and B(59)) xor (A(112) and B(58)) xor (A(113) and B(57)) xor (A(114) and B(56)) xor (A(115) and B(55)) xor (A(116) and B(54)) xor (A(117) and B(53)) xor (A(118) and B(52)) xor (A(119) and B(51)) xor (A(120) and B(50)) xor (A(121) and B(49)) xor (A(122) and B(48)) xor (A(123) and B(47)) xor (A(124) and B(46)) xor (A(125) and B(45)) xor (A(126) and B(44)) xor (A(48) and B(127)) xor (A(49) and B(126)) xor (A(50) and B(125)) xor (A(51) and B(124)) xor (A(52) and B(123)) xor (A(53) and B(122)) xor (A(54) and B(121)) xor (A(55) and B(120)) xor (A(56) and B(119)) xor (A(57) and B(118)) xor (A(58) and B(117)) xor (A(59) and B(116)) xor (A(60) and B(115)) xor (A(61) and B(114)) xor (A(62) and B(113)) xor (A(63) and B(112)) xor (A(64) and B(111)) xor (A(65) and B(110)) xor (A(66) and B(109)) xor (A(67) and B(108)) xor (A(68) and B(107)) xor (A(69) and B(106)) xor (A(70) and B(105)) xor (A(71) and B(104)) xor (A(72) and B(103)) xor (A(73) and B(102)) xor (A(74) and B(101)) xor (A(75) and B(100)) xor (A(76) and B(99)) xor (A(77) and B(98)) xor (A(78) and B(97)) xor (A(79) and B(96)) xor (A(80) and B(95)) xor (A(81) and B(94)) xor (A(82) and B(93)) xor (A(83) and B(92)) xor (A(84) and B(91)) xor (A(85) and B(90)) xor (A(86) and B(89)) xor (A(87) and B(88)) xor (A(88) and B(87)) xor (A(89) and B(86)) xor (A(90) and B(85)) xor (A(91) and B(84)) xor (A(92) and B(83)) xor (A(93) and B(82)) xor (A(94) and B(81)) xor (A(95) and B(80)) xor (A(96) and B(79)) xor (A(97) and B(78)) xor (A(98) and B(77)) xor (A(99) and B(76)) xor (A(100) and B(75)) xor (A(101) and B(74)) xor (A(102) and B(73)) xor (A(103) and B(72)) xor (A(104) and B(71)) xor (A(105) and B(70)) xor (A(106) and B(69)) xor (A(107) and B(68)) xor (A(108) and B(67)) xor (A(109) and B(66)) xor (A(110) and B(65)) xor (A(111) and B(64)) xor (A(112) and B(63)) xor (A(113) and B(62)) xor (A(114) and B(61)) xor (A(115) and B(60)) xor (A(116) and B(59)) xor (A(117) and B(58)) xor (A(118) and B(57)) xor (A(119) and B(56)) xor (A(120) and B(55)) xor (A(121) and B(54)) xor (A(122) and B(53)) xor (A(123) and B(52)) xor (A(124) and B(51)) xor (A(125) and B(50)) xor (A(126) and B(49)) xor (A(49) and B(127)) xor (A(50) and B(126)) xor (A(51) and B(125)) xor (A(52) and B(124)) xor (A(53) and B(123)) xor (A(54) and B(122)) xor (A(55) and B(121)) xor (A(56) and B(120)) xor (A(57) and B(119)) xor (A(58) and B(118)) xor (A(59) and B(117)) xor (A(60) and B(116)) xor (A(61) and B(115)) xor (A(62) and B(114)) xor (A(63) and B(113)) xor (A(64) and B(112)) xor (A(65) and B(111)) xor (A(66) and B(110)) xor (A(67) and B(109)) xor (A(68) and B(108)) xor (A(69) and B(107)) xor (A(70) and B(106)) xor (A(71) and B(105)) xor (A(72) and B(104)) xor (A(73) and B(103)) xor (A(74) and B(102)) xor (A(75) and B(101)) xor (A(76) and B(100)) xor (A(77) and B(99)) xor (A(78) and B(98)) xor (A(79) and B(97)) xor (A(80) and B(96)) xor (A(81) and B(95)) xor (A(82) and B(94)) xor (A(83) and B(93)) xor (A(84) and B(92)) xor (A(85) and B(91)) xor (A(86) and B(90)) xor (A(87) and B(89)) xor (A(88) and B(88)) xor (A(89) and B(87)) xor (A(90) and B(86)) xor (A(91) and B(85)) xor (A(92) and B(84)) xor (A(93) and B(83)) xor (A(94) and B(82)) xor (A(95) and B(81)) xor (A(96) and B(80)) xor (A(97) and B(79)) xor (A(98) and B(78)) xor (A(99) and B(77)) xor (A(100) and B(76)) xor (A(101) and B(75)) xor (A(102) and B(74)) xor (A(103) and B(73)) xor (A(104) and B(72)) xor (A(105) and B(71)) xor (A(106) and B(70)) xor (A(107) and B(69)) xor (A(108) and B(68)) xor (A(109) and B(67)) xor (A(110) and B(66)) xor (A(111) and B(65)) xor (A(112) and B(64)) xor (A(113) and B(63)) xor (A(114) and B(62)) xor (A(115) and B(61)) xor (A(116) and B(60)) xor (A(117) and B(59)) xor (A(118) and B(58)) xor (A(119) and B(57)) xor (A(120) and B(56)) xor (A(121) and B(55)) xor (A(122) and B(54)) xor (A(123) and B(53)) xor (A(124) and B(52)) xor (A(125) and B(51)) xor (A(126) and B(50)) xor (A(50) and B(127)) xor (A(51) and B(126)) xor (A(52) and B(125)) xor (A(53) and B(124)) xor (A(54) and B(123)) xor (A(55) and B(122)) xor (A(56) and B(121)) xor (A(57) and B(120)) xor (A(58) and B(119)) xor (A(59) and B(118)) xor (A(60) and B(117)) xor (A(61) and B(116)) xor (A(62) and B(115)) xor (A(63) and B(114)) xor (A(64) and B(113)) xor (A(65) and B(112)) xor (A(66) and B(111)) xor (A(67) and B(110)) xor (A(68) and B(109)) xor (A(69) and B(108)) xor (A(70) and B(107)) xor (A(71) and B(106)) xor (A(72) and B(105)) xor (A(73) and B(104)) xor (A(74) and B(103)) xor (A(75) and B(102)) xor (A(76) and B(101)) xor (A(77) and B(100)) xor (A(78) and B(99)) xor (A(79) and B(98)) xor (A(80) and B(97)) xor (A(81) and B(96)) xor (A(82) and B(95)) xor (A(83) and B(94)) xor (A(84) and B(93)) xor (A(85) and B(92)) xor (A(86) and B(91)) xor (A(87) and B(90)) xor (A(88) and B(89)) xor (A(89) and B(88)) xor (A(90) and B(87)) xor (A(91) and B(86)) xor (A(92) and B(85)) xor (A(93) and B(84)) xor (A(94) and B(83)) xor (A(95) and B(82)) xor (A(96) and B(81)) xor (A(97) and B(80)) xor (A(98) and B(79)) xor (A(99) and B(78)) xor (A(100) and B(77)) xor (A(101) and B(76)) xor (A(102) and B(75)) xor (A(103) and B(74)) xor (A(104) and B(73)) xor (A(105) and B(72)) xor (A(106) and B(71)) xor (A(107) and B(70)) xor (A(108) and B(69)) xor (A(109) and B(68)) xor (A(110) and B(67)) xor (A(111) and B(66)) xor (A(112) and B(65)) xor (A(113) and B(64)) xor (A(114) and B(63)) xor (A(115) and B(62)) xor (A(116) and B(61)) xor (A(117) and B(60)) xor (A(118) and B(59)) xor (A(119) and B(58)) xor (A(120) and B(57)) xor (A(121) and B(56)) xor (A(122) and B(55)) xor (A(123) and B(54)) xor (A(124) and B(53)) xor (A(125) and B(52)) xor (A(126) and B(52));
    C(51)  <= (A(0) and B(51)) xor (A(1) and B(50)) xor (A(2) and B(49)) xor (A(3) and B(48)) xor (A(4) and B(47)) xor (A(5) and B(46)) xor (A(6) and B(45)) xor (A(7) and B(44)) xor (A(8) and B(43)) xor (A(9) and B(42)) xor (A(10) and B(41)) xor (A(11) and B(40)) xor (A(12) and B(39)) xor (A(13) and B(38)) xor (A(14) and B(37)) xor (A(15) and B(36)) xor (A(16) and B(35)) xor (A(17) and B(34)) xor (A(18) and B(33)) xor (A(19) and B(32)) xor (A(20) and B(31)) xor (A(21) and B(30)) xor (A(23) and B(29)) xor (A(23) and B(28)) xor (A(24) and B(27)) xor (A(25) and B(26)) xor (A(26) and B(25)) xor (A(27) and B(24)) xor (A(28) and B(23)) xor (A(29) and B(23)) xor (A(30) and B(21)) xor (A(31) and B(20)) xor (A(32) and B(19)) xor (A(33) and B(18)) xor (A(34) and B(17)) xor (A(35) and B(16)) xor (A(36) and B(15)) xor (A(37) and B(14)) xor (A(38) and B(13)) xor (A(39) and B(12)) xor (A(40) and B(11)) xor (A(41) and B(10)) xor (A(42) and B(9)) xor (A(43) and B(8)) xor (A(44) and B(7)) xor (A(45) and B(6)) xor (A(46) and B(5)) xor (A(47) and B(4)) xor (A(48) and B(3)) xor (A(49) and B(2)) xor (A(50) and B(1)) xor (A(51) and B(0)) xor (A(44) and B(127)) xor (A(45) and B(126)) xor (A(46) and B(125)) xor (A(47) and B(124)) xor (A(48) and B(123)) xor (A(49) and B(122)) xor (A(50) and B(121)) xor (A(51) and B(120)) xor (A(52) and B(119)) xor (A(53) and B(118)) xor (A(54) and B(117)) xor (A(55) and B(116)) xor (A(56) and B(115)) xor (A(57) and B(114)) xor (A(58) and B(113)) xor (A(59) and B(112)) xor (A(60) and B(111)) xor (A(61) and B(110)) xor (A(62) and B(109)) xor (A(63) and B(108)) xor (A(64) and B(107)) xor (A(65) and B(106)) xor (A(66) and B(105)) xor (A(67) and B(104)) xor (A(68) and B(103)) xor (A(69) and B(102)) xor (A(70) and B(101)) xor (A(71) and B(100)) xor (A(72) and B(99)) xor (A(73) and B(98)) xor (A(74) and B(97)) xor (A(75) and B(96)) xor (A(76) and B(95)) xor (A(77) and B(94)) xor (A(78) and B(93)) xor (A(79) and B(92)) xor (A(80) and B(91)) xor (A(81) and B(90)) xor (A(82) and B(89)) xor (A(83) and B(88)) xor (A(84) and B(87)) xor (A(85) and B(86)) xor (A(86) and B(85)) xor (A(87) and B(84)) xor (A(88) and B(83)) xor (A(89) and B(82)) xor (A(90) and B(81)) xor (A(91) and B(80)) xor (A(92) and B(79)) xor (A(93) and B(78)) xor (A(94) and B(77)) xor (A(95) and B(76)) xor (A(96) and B(75)) xor (A(97) and B(74)) xor (A(98) and B(73)) xor (A(99) and B(72)) xor (A(100) and B(71)) xor (A(101) and B(70)) xor (A(102) and B(69)) xor (A(103) and B(68)) xor (A(104) and B(67)) xor (A(105) and B(66)) xor (A(106) and B(65)) xor (A(107) and B(64)) xor (A(108) and B(63)) xor (A(109) and B(62)) xor (A(110) and B(61)) xor (A(111) and B(60)) xor (A(112) and B(59)) xor (A(113) and B(58)) xor (A(114) and B(57)) xor (A(115) and B(56)) xor (A(116) and B(55)) xor (A(117) and B(54)) xor (A(118) and B(53)) xor (A(119) and B(52)) xor (A(120) and B(51)) xor (A(121) and B(50)) xor (A(122) and B(49)) xor (A(123) and B(48)) xor (A(124) and B(47)) xor (A(125) and B(46)) xor (A(126) and B(45)) xor (A(49) and B(127)) xor (A(50) and B(126)) xor (A(51) and B(125)) xor (A(52) and B(124)) xor (A(53) and B(123)) xor (A(54) and B(122)) xor (A(55) and B(121)) xor (A(56) and B(120)) xor (A(57) and B(119)) xor (A(58) and B(118)) xor (A(59) and B(117)) xor (A(60) and B(116)) xor (A(61) and B(115)) xor (A(62) and B(114)) xor (A(63) and B(113)) xor (A(64) and B(112)) xor (A(65) and B(111)) xor (A(66) and B(110)) xor (A(67) and B(109)) xor (A(68) and B(108)) xor (A(69) and B(107)) xor (A(70) and B(106)) xor (A(71) and B(105)) xor (A(72) and B(104)) xor (A(73) and B(103)) xor (A(74) and B(102)) xor (A(75) and B(101)) xor (A(76) and B(100)) xor (A(77) and B(99)) xor (A(78) and B(98)) xor (A(79) and B(97)) xor (A(80) and B(96)) xor (A(81) and B(95)) xor (A(82) and B(94)) xor (A(83) and B(93)) xor (A(84) and B(92)) xor (A(85) and B(91)) xor (A(86) and B(90)) xor (A(87) and B(89)) xor (A(88) and B(88)) xor (A(89) and B(87)) xor (A(90) and B(86)) xor (A(91) and B(85)) xor (A(92) and B(84)) xor (A(93) and B(83)) xor (A(94) and B(82)) xor (A(95) and B(81)) xor (A(96) and B(80)) xor (A(97) and B(79)) xor (A(98) and B(78)) xor (A(99) and B(77)) xor (A(100) and B(76)) xor (A(101) and B(75)) xor (A(102) and B(74)) xor (A(103) and B(73)) xor (A(104) and B(72)) xor (A(105) and B(71)) xor (A(106) and B(70)) xor (A(107) and B(69)) xor (A(108) and B(68)) xor (A(109) and B(67)) xor (A(110) and B(66)) xor (A(111) and B(65)) xor (A(112) and B(64)) xor (A(113) and B(63)) xor (A(114) and B(62)) xor (A(115) and B(61)) xor (A(116) and B(60)) xor (A(117) and B(59)) xor (A(118) and B(58)) xor (A(119) and B(57)) xor (A(120) and B(56)) xor (A(121) and B(55)) xor (A(122) and B(54)) xor (A(123) and B(53)) xor (A(124) and B(52)) xor (A(125) and B(51)) xor (A(126) and B(50)) xor (A(50) and B(127)) xor (A(51) and B(126)) xor (A(52) and B(125)) xor (A(53) and B(124)) xor (A(54) and B(123)) xor (A(55) and B(122)) xor (A(56) and B(121)) xor (A(57) and B(120)) xor (A(58) and B(119)) xor (A(59) and B(118)) xor (A(60) and B(117)) xor (A(61) and B(116)) xor (A(62) and B(115)) xor (A(63) and B(114)) xor (A(64) and B(113)) xor (A(65) and B(112)) xor (A(66) and B(111)) xor (A(67) and B(110)) xor (A(68) and B(109)) xor (A(69) and B(108)) xor (A(70) and B(107)) xor (A(71) and B(106)) xor (A(72) and B(105)) xor (A(73) and B(104)) xor (A(74) and B(103)) xor (A(75) and B(102)) xor (A(76) and B(101)) xor (A(77) and B(100)) xor (A(78) and B(99)) xor (A(79) and B(98)) xor (A(80) and B(97)) xor (A(81) and B(96)) xor (A(82) and B(95)) xor (A(83) and B(94)) xor (A(84) and B(93)) xor (A(85) and B(92)) xor (A(86) and B(91)) xor (A(87) and B(90)) xor (A(88) and B(89)) xor (A(89) and B(88)) xor (A(90) and B(87)) xor (A(91) and B(86)) xor (A(92) and B(85)) xor (A(93) and B(84)) xor (A(94) and B(83)) xor (A(95) and B(82)) xor (A(96) and B(81)) xor (A(97) and B(80)) xor (A(98) and B(79)) xor (A(99) and B(78)) xor (A(100) and B(77)) xor (A(101) and B(76)) xor (A(102) and B(75)) xor (A(103) and B(74)) xor (A(104) and B(73)) xor (A(105) and B(72)) xor (A(106) and B(71)) xor (A(107) and B(70)) xor (A(108) and B(69)) xor (A(109) and B(68)) xor (A(110) and B(67)) xor (A(111) and B(66)) xor (A(112) and B(65)) xor (A(113) and B(64)) xor (A(114) and B(63)) xor (A(115) and B(62)) xor (A(116) and B(61)) xor (A(117) and B(60)) xor (A(118) and B(59)) xor (A(119) and B(58)) xor (A(120) and B(57)) xor (A(121) and B(56)) xor (A(122) and B(55)) xor (A(123) and B(54)) xor (A(124) and B(53)) xor (A(125) and B(52)) xor (A(126) and B(51)) xor (A(51) and B(127)) xor (A(52) and B(126)) xor (A(53) and B(125)) xor (A(54) and B(124)) xor (A(55) and B(123)) xor (A(56) and B(122)) xor (A(57) and B(121)) xor (A(58) and B(120)) xor (A(59) and B(119)) xor (A(60) and B(118)) xor (A(61) and B(117)) xor (A(62) and B(116)) xor (A(63) and B(115)) xor (A(64) and B(114)) xor (A(65) and B(113)) xor (A(66) and B(112)) xor (A(67) and B(111)) xor (A(68) and B(110)) xor (A(69) and B(109)) xor (A(70) and B(108)) xor (A(71) and B(107)) xor (A(72) and B(106)) xor (A(73) and B(105)) xor (A(74) and B(104)) xor (A(75) and B(103)) xor (A(76) and B(102)) xor (A(77) and B(101)) xor (A(78) and B(100)) xor (A(79) and B(99)) xor (A(80) and B(98)) xor (A(81) and B(97)) xor (A(82) and B(96)) xor (A(83) and B(95)) xor (A(84) and B(94)) xor (A(85) and B(93)) xor (A(86) and B(92)) xor (A(87) and B(91)) xor (A(88) and B(90)) xor (A(89) and B(89)) xor (A(90) and B(88)) xor (A(91) and B(87)) xor (A(92) and B(86)) xor (A(93) and B(85)) xor (A(94) and B(84)) xor (A(95) and B(83)) xor (A(96) and B(82)) xor (A(97) and B(81)) xor (A(98) and B(80)) xor (A(99) and B(79)) xor (A(100) and B(78)) xor (A(101) and B(77)) xor (A(102) and B(76)) xor (A(103) and B(75)) xor (A(104) and B(74)) xor (A(105) and B(73)) xor (A(106) and B(72)) xor (A(107) and B(71)) xor (A(108) and B(70)) xor (A(109) and B(69)) xor (A(110) and B(68)) xor (A(111) and B(67)) xor (A(112) and B(66)) xor (A(113) and B(65)) xor (A(114) and B(64)) xor (A(115) and B(63)) xor (A(116) and B(62)) xor (A(117) and B(61)) xor (A(118) and B(60)) xor (A(119) and B(59)) xor (A(120) and B(58)) xor (A(121) and B(57)) xor (A(122) and B(56)) xor (A(123) and B(55)) xor (A(124) and B(54)) xor (A(125) and B(53)) xor (A(126) and B(53));
    C(52)  <= (A(0) and B(52)) xor (A(1) and B(51)) xor (A(2) and B(50)) xor (A(3) and B(49)) xor (A(4) and B(48)) xor (A(5) and B(47)) xor (A(6) and B(46)) xor (A(7) and B(45)) xor (A(8) and B(44)) xor (A(9) and B(43)) xor (A(10) and B(42)) xor (A(11) and B(41)) xor (A(12) and B(40)) xor (A(13) and B(39)) xor (A(14) and B(38)) xor (A(15) and B(37)) xor (A(16) and B(36)) xor (A(17) and B(35)) xor (A(18) and B(34)) xor (A(19) and B(33)) xor (A(20) and B(32)) xor (A(21) and B(31)) xor (A(23) and B(30)) xor (A(23) and B(29)) xor (A(24) and B(28)) xor (A(25) and B(27)) xor (A(26) and B(26)) xor (A(27) and B(25)) xor (A(28) and B(24)) xor (A(29) and B(23)) xor (A(30) and B(23)) xor (A(31) and B(21)) xor (A(32) and B(20)) xor (A(33) and B(19)) xor (A(34) and B(18)) xor (A(35) and B(17)) xor (A(36) and B(16)) xor (A(37) and B(15)) xor (A(38) and B(14)) xor (A(39) and B(13)) xor (A(40) and B(12)) xor (A(41) and B(11)) xor (A(42) and B(10)) xor (A(43) and B(9)) xor (A(44) and B(8)) xor (A(45) and B(7)) xor (A(46) and B(6)) xor (A(47) and B(5)) xor (A(48) and B(4)) xor (A(49) and B(3)) xor (A(50) and B(2)) xor (A(51) and B(1)) xor (A(52) and B(0)) xor (A(45) and B(127)) xor (A(46) and B(126)) xor (A(47) and B(125)) xor (A(48) and B(124)) xor (A(49) and B(123)) xor (A(50) and B(122)) xor (A(51) and B(121)) xor (A(52) and B(120)) xor (A(53) and B(119)) xor (A(54) and B(118)) xor (A(55) and B(117)) xor (A(56) and B(116)) xor (A(57) and B(115)) xor (A(58) and B(114)) xor (A(59) and B(113)) xor (A(60) and B(112)) xor (A(61) and B(111)) xor (A(62) and B(110)) xor (A(63) and B(109)) xor (A(64) and B(108)) xor (A(65) and B(107)) xor (A(66) and B(106)) xor (A(67) and B(105)) xor (A(68) and B(104)) xor (A(69) and B(103)) xor (A(70) and B(102)) xor (A(71) and B(101)) xor (A(72) and B(100)) xor (A(73) and B(99)) xor (A(74) and B(98)) xor (A(75) and B(97)) xor (A(76) and B(96)) xor (A(77) and B(95)) xor (A(78) and B(94)) xor (A(79) and B(93)) xor (A(80) and B(92)) xor (A(81) and B(91)) xor (A(82) and B(90)) xor (A(83) and B(89)) xor (A(84) and B(88)) xor (A(85) and B(87)) xor (A(86) and B(86)) xor (A(87) and B(85)) xor (A(88) and B(84)) xor (A(89) and B(83)) xor (A(90) and B(82)) xor (A(91) and B(81)) xor (A(92) and B(80)) xor (A(93) and B(79)) xor (A(94) and B(78)) xor (A(95) and B(77)) xor (A(96) and B(76)) xor (A(97) and B(75)) xor (A(98) and B(74)) xor (A(99) and B(73)) xor (A(100) and B(72)) xor (A(101) and B(71)) xor (A(102) and B(70)) xor (A(103) and B(69)) xor (A(104) and B(68)) xor (A(105) and B(67)) xor (A(106) and B(66)) xor (A(107) and B(65)) xor (A(108) and B(64)) xor (A(109) and B(63)) xor (A(110) and B(62)) xor (A(111) and B(61)) xor (A(112) and B(60)) xor (A(113) and B(59)) xor (A(114) and B(58)) xor (A(115) and B(57)) xor (A(116) and B(56)) xor (A(117) and B(55)) xor (A(118) and B(54)) xor (A(119) and B(53)) xor (A(120) and B(52)) xor (A(121) and B(51)) xor (A(122) and B(50)) xor (A(123) and B(49)) xor (A(124) and B(48)) xor (A(125) and B(47)) xor (A(126) and B(46)) xor (A(50) and B(127)) xor (A(51) and B(126)) xor (A(52) and B(125)) xor (A(53) and B(124)) xor (A(54) and B(123)) xor (A(55) and B(122)) xor (A(56) and B(121)) xor (A(57) and B(120)) xor (A(58) and B(119)) xor (A(59) and B(118)) xor (A(60) and B(117)) xor (A(61) and B(116)) xor (A(62) and B(115)) xor (A(63) and B(114)) xor (A(64) and B(113)) xor (A(65) and B(112)) xor (A(66) and B(111)) xor (A(67) and B(110)) xor (A(68) and B(109)) xor (A(69) and B(108)) xor (A(70) and B(107)) xor (A(71) and B(106)) xor (A(72) and B(105)) xor (A(73) and B(104)) xor (A(74) and B(103)) xor (A(75) and B(102)) xor (A(76) and B(101)) xor (A(77) and B(100)) xor (A(78) and B(99)) xor (A(79) and B(98)) xor (A(80) and B(97)) xor (A(81) and B(96)) xor (A(82) and B(95)) xor (A(83) and B(94)) xor (A(84) and B(93)) xor (A(85) and B(92)) xor (A(86) and B(91)) xor (A(87) and B(90)) xor (A(88) and B(89)) xor (A(89) and B(88)) xor (A(90) and B(87)) xor (A(91) and B(86)) xor (A(92) and B(85)) xor (A(93) and B(84)) xor (A(94) and B(83)) xor (A(95) and B(82)) xor (A(96) and B(81)) xor (A(97) and B(80)) xor (A(98) and B(79)) xor (A(99) and B(78)) xor (A(100) and B(77)) xor (A(101) and B(76)) xor (A(102) and B(75)) xor (A(103) and B(74)) xor (A(104) and B(73)) xor (A(105) and B(72)) xor (A(106) and B(71)) xor (A(107) and B(70)) xor (A(108) and B(69)) xor (A(109) and B(68)) xor (A(110) and B(67)) xor (A(111) and B(66)) xor (A(112) and B(65)) xor (A(113) and B(64)) xor (A(114) and B(63)) xor (A(115) and B(62)) xor (A(116) and B(61)) xor (A(117) and B(60)) xor (A(118) and B(59)) xor (A(119) and B(58)) xor (A(120) and B(57)) xor (A(121) and B(56)) xor (A(122) and B(55)) xor (A(123) and B(54)) xor (A(124) and B(53)) xor (A(125) and B(52)) xor (A(126) and B(51)) xor (A(51) and B(127)) xor (A(52) and B(126)) xor (A(53) and B(125)) xor (A(54) and B(124)) xor (A(55) and B(123)) xor (A(56) and B(122)) xor (A(57) and B(121)) xor (A(58) and B(120)) xor (A(59) and B(119)) xor (A(60) and B(118)) xor (A(61) and B(117)) xor (A(62) and B(116)) xor (A(63) and B(115)) xor (A(64) and B(114)) xor (A(65) and B(113)) xor (A(66) and B(112)) xor (A(67) and B(111)) xor (A(68) and B(110)) xor (A(69) and B(109)) xor (A(70) and B(108)) xor (A(71) and B(107)) xor (A(72) and B(106)) xor (A(73) and B(105)) xor (A(74) and B(104)) xor (A(75) and B(103)) xor (A(76) and B(102)) xor (A(77) and B(101)) xor (A(78) and B(100)) xor (A(79) and B(99)) xor (A(80) and B(98)) xor (A(81) and B(97)) xor (A(82) and B(96)) xor (A(83) and B(95)) xor (A(84) and B(94)) xor (A(85) and B(93)) xor (A(86) and B(92)) xor (A(87) and B(91)) xor (A(88) and B(90)) xor (A(89) and B(89)) xor (A(90) and B(88)) xor (A(91) and B(87)) xor (A(92) and B(86)) xor (A(93) and B(85)) xor (A(94) and B(84)) xor (A(95) and B(83)) xor (A(96) and B(82)) xor (A(97) and B(81)) xor (A(98) and B(80)) xor (A(99) and B(79)) xor (A(100) and B(78)) xor (A(101) and B(77)) xor (A(102) and B(76)) xor (A(103) and B(75)) xor (A(104) and B(74)) xor (A(105) and B(73)) xor (A(106) and B(72)) xor (A(107) and B(71)) xor (A(108) and B(70)) xor (A(109) and B(69)) xor (A(110) and B(68)) xor (A(111) and B(67)) xor (A(112) and B(66)) xor (A(113) and B(65)) xor (A(114) and B(64)) xor (A(115) and B(63)) xor (A(116) and B(62)) xor (A(117) and B(61)) xor (A(118) and B(60)) xor (A(119) and B(59)) xor (A(120) and B(58)) xor (A(121) and B(57)) xor (A(122) and B(56)) xor (A(123) and B(55)) xor (A(124) and B(54)) xor (A(125) and B(53)) xor (A(126) and B(52)) xor (A(52) and B(127)) xor (A(53) and B(126)) xor (A(54) and B(125)) xor (A(55) and B(124)) xor (A(56) and B(123)) xor (A(57) and B(122)) xor (A(58) and B(121)) xor (A(59) and B(120)) xor (A(60) and B(119)) xor (A(61) and B(118)) xor (A(62) and B(117)) xor (A(63) and B(116)) xor (A(64) and B(115)) xor (A(65) and B(114)) xor (A(66) and B(113)) xor (A(67) and B(112)) xor (A(68) and B(111)) xor (A(69) and B(110)) xor (A(70) and B(109)) xor (A(71) and B(108)) xor (A(72) and B(107)) xor (A(73) and B(106)) xor (A(74) and B(105)) xor (A(75) and B(104)) xor (A(76) and B(103)) xor (A(77) and B(102)) xor (A(78) and B(101)) xor (A(79) and B(100)) xor (A(80) and B(99)) xor (A(81) and B(98)) xor (A(82) and B(97)) xor (A(83) and B(96)) xor (A(84) and B(95)) xor (A(85) and B(94)) xor (A(86) and B(93)) xor (A(87) and B(92)) xor (A(88) and B(91)) xor (A(89) and B(90)) xor (A(90) and B(89)) xor (A(91) and B(88)) xor (A(92) and B(87)) xor (A(93) and B(86)) xor (A(94) and B(85)) xor (A(95) and B(84)) xor (A(96) and B(83)) xor (A(97) and B(82)) xor (A(98) and B(81)) xor (A(99) and B(80)) xor (A(100) and B(79)) xor (A(101) and B(78)) xor (A(102) and B(77)) xor (A(103) and B(76)) xor (A(104) and B(75)) xor (A(105) and B(74)) xor (A(106) and B(73)) xor (A(107) and B(72)) xor (A(108) and B(71)) xor (A(109) and B(70)) xor (A(110) and B(69)) xor (A(111) and B(68)) xor (A(112) and B(67)) xor (A(113) and B(66)) xor (A(114) and B(65)) xor (A(115) and B(64)) xor (A(116) and B(63)) xor (A(117) and B(62)) xor (A(118) and B(61)) xor (A(119) and B(60)) xor (A(120) and B(59)) xor (A(121) and B(58)) xor (A(122) and B(57)) xor (A(123) and B(56)) xor (A(124) and B(55)) xor (A(125) and B(54)) xor (A(126) and B(54));
    C(53)  <= (A(0) and B(53)) xor (A(1) and B(52)) xor (A(2) and B(51)) xor (A(3) and B(50)) xor (A(4) and B(49)) xor (A(5) and B(48)) xor (A(6) and B(47)) xor (A(7) and B(46)) xor (A(8) and B(45)) xor (A(9) and B(44)) xor (A(10) and B(43)) xor (A(11) and B(42)) xor (A(12) and B(41)) xor (A(13) and B(40)) xor (A(14) and B(39)) xor (A(15) and B(38)) xor (A(16) and B(37)) xor (A(17) and B(36)) xor (A(18) and B(35)) xor (A(19) and B(34)) xor (A(20) and B(33)) xor (A(21) and B(32)) xor (A(23) and B(31)) xor (A(23) and B(30)) xor (A(24) and B(29)) xor (A(25) and B(28)) xor (A(26) and B(27)) xor (A(27) and B(26)) xor (A(28) and B(25)) xor (A(29) and B(24)) xor (A(30) and B(23)) xor (A(31) and B(23)) xor (A(32) and B(21)) xor (A(33) and B(20)) xor (A(34) and B(19)) xor (A(35) and B(18)) xor (A(36) and B(17)) xor (A(37) and B(16)) xor (A(38) and B(15)) xor (A(39) and B(14)) xor (A(40) and B(13)) xor (A(41) and B(12)) xor (A(42) and B(11)) xor (A(43) and B(10)) xor (A(44) and B(9)) xor (A(45) and B(8)) xor (A(46) and B(7)) xor (A(47) and B(6)) xor (A(48) and B(5)) xor (A(49) and B(4)) xor (A(50) and B(3)) xor (A(51) and B(2)) xor (A(52) and B(1)) xor (A(53) and B(0)) xor (A(46) and B(127)) xor (A(47) and B(126)) xor (A(48) and B(125)) xor (A(49) and B(124)) xor (A(50) and B(123)) xor (A(51) and B(122)) xor (A(52) and B(121)) xor (A(53) and B(120)) xor (A(54) and B(119)) xor (A(55) and B(118)) xor (A(56) and B(117)) xor (A(57) and B(116)) xor (A(58) and B(115)) xor (A(59) and B(114)) xor (A(60) and B(113)) xor (A(61) and B(112)) xor (A(62) and B(111)) xor (A(63) and B(110)) xor (A(64) and B(109)) xor (A(65) and B(108)) xor (A(66) and B(107)) xor (A(67) and B(106)) xor (A(68) and B(105)) xor (A(69) and B(104)) xor (A(70) and B(103)) xor (A(71) and B(102)) xor (A(72) and B(101)) xor (A(73) and B(100)) xor (A(74) and B(99)) xor (A(75) and B(98)) xor (A(76) and B(97)) xor (A(77) and B(96)) xor (A(78) and B(95)) xor (A(79) and B(94)) xor (A(80) and B(93)) xor (A(81) and B(92)) xor (A(82) and B(91)) xor (A(83) and B(90)) xor (A(84) and B(89)) xor (A(85) and B(88)) xor (A(86) and B(87)) xor (A(87) and B(86)) xor (A(88) and B(85)) xor (A(89) and B(84)) xor (A(90) and B(83)) xor (A(91) and B(82)) xor (A(92) and B(81)) xor (A(93) and B(80)) xor (A(94) and B(79)) xor (A(95) and B(78)) xor (A(96) and B(77)) xor (A(97) and B(76)) xor (A(98) and B(75)) xor (A(99) and B(74)) xor (A(100) and B(73)) xor (A(101) and B(72)) xor (A(102) and B(71)) xor (A(103) and B(70)) xor (A(104) and B(69)) xor (A(105) and B(68)) xor (A(106) and B(67)) xor (A(107) and B(66)) xor (A(108) and B(65)) xor (A(109) and B(64)) xor (A(110) and B(63)) xor (A(111) and B(62)) xor (A(112) and B(61)) xor (A(113) and B(60)) xor (A(114) and B(59)) xor (A(115) and B(58)) xor (A(116) and B(57)) xor (A(117) and B(56)) xor (A(118) and B(55)) xor (A(119) and B(54)) xor (A(120) and B(53)) xor (A(121) and B(52)) xor (A(122) and B(51)) xor (A(123) and B(50)) xor (A(124) and B(49)) xor (A(125) and B(48)) xor (A(126) and B(47)) xor (A(51) and B(127)) xor (A(52) and B(126)) xor (A(53) and B(125)) xor (A(54) and B(124)) xor (A(55) and B(123)) xor (A(56) and B(122)) xor (A(57) and B(121)) xor (A(58) and B(120)) xor (A(59) and B(119)) xor (A(60) and B(118)) xor (A(61) and B(117)) xor (A(62) and B(116)) xor (A(63) and B(115)) xor (A(64) and B(114)) xor (A(65) and B(113)) xor (A(66) and B(112)) xor (A(67) and B(111)) xor (A(68) and B(110)) xor (A(69) and B(109)) xor (A(70) and B(108)) xor (A(71) and B(107)) xor (A(72) and B(106)) xor (A(73) and B(105)) xor (A(74) and B(104)) xor (A(75) and B(103)) xor (A(76) and B(102)) xor (A(77) and B(101)) xor (A(78) and B(100)) xor (A(79) and B(99)) xor (A(80) and B(98)) xor (A(81) and B(97)) xor (A(82) and B(96)) xor (A(83) and B(95)) xor (A(84) and B(94)) xor (A(85) and B(93)) xor (A(86) and B(92)) xor (A(87) and B(91)) xor (A(88) and B(90)) xor (A(89) and B(89)) xor (A(90) and B(88)) xor (A(91) and B(87)) xor (A(92) and B(86)) xor (A(93) and B(85)) xor (A(94) and B(84)) xor (A(95) and B(83)) xor (A(96) and B(82)) xor (A(97) and B(81)) xor (A(98) and B(80)) xor (A(99) and B(79)) xor (A(100) and B(78)) xor (A(101) and B(77)) xor (A(102) and B(76)) xor (A(103) and B(75)) xor (A(104) and B(74)) xor (A(105) and B(73)) xor (A(106) and B(72)) xor (A(107) and B(71)) xor (A(108) and B(70)) xor (A(109) and B(69)) xor (A(110) and B(68)) xor (A(111) and B(67)) xor (A(112) and B(66)) xor (A(113) and B(65)) xor (A(114) and B(64)) xor (A(115) and B(63)) xor (A(116) and B(62)) xor (A(117) and B(61)) xor (A(118) and B(60)) xor (A(119) and B(59)) xor (A(120) and B(58)) xor (A(121) and B(57)) xor (A(122) and B(56)) xor (A(123) and B(55)) xor (A(124) and B(54)) xor (A(125) and B(53)) xor (A(126) and B(52)) xor (A(52) and B(127)) xor (A(53) and B(126)) xor (A(54) and B(125)) xor (A(55) and B(124)) xor (A(56) and B(123)) xor (A(57) and B(122)) xor (A(58) and B(121)) xor (A(59) and B(120)) xor (A(60) and B(119)) xor (A(61) and B(118)) xor (A(62) and B(117)) xor (A(63) and B(116)) xor (A(64) and B(115)) xor (A(65) and B(114)) xor (A(66) and B(113)) xor (A(67) and B(112)) xor (A(68) and B(111)) xor (A(69) and B(110)) xor (A(70) and B(109)) xor (A(71) and B(108)) xor (A(72) and B(107)) xor (A(73) and B(106)) xor (A(74) and B(105)) xor (A(75) and B(104)) xor (A(76) and B(103)) xor (A(77) and B(102)) xor (A(78) and B(101)) xor (A(79) and B(100)) xor (A(80) and B(99)) xor (A(81) and B(98)) xor (A(82) and B(97)) xor (A(83) and B(96)) xor (A(84) and B(95)) xor (A(85) and B(94)) xor (A(86) and B(93)) xor (A(87) and B(92)) xor (A(88) and B(91)) xor (A(89) and B(90)) xor (A(90) and B(89)) xor (A(91) and B(88)) xor (A(92) and B(87)) xor (A(93) and B(86)) xor (A(94) and B(85)) xor (A(95) and B(84)) xor (A(96) and B(83)) xor (A(97) and B(82)) xor (A(98) and B(81)) xor (A(99) and B(80)) xor (A(100) and B(79)) xor (A(101) and B(78)) xor (A(102) and B(77)) xor (A(103) and B(76)) xor (A(104) and B(75)) xor (A(105) and B(74)) xor (A(106) and B(73)) xor (A(107) and B(72)) xor (A(108) and B(71)) xor (A(109) and B(70)) xor (A(110) and B(69)) xor (A(111) and B(68)) xor (A(112) and B(67)) xor (A(113) and B(66)) xor (A(114) and B(65)) xor (A(115) and B(64)) xor (A(116) and B(63)) xor (A(117) and B(62)) xor (A(118) and B(61)) xor (A(119) and B(60)) xor (A(120) and B(59)) xor (A(121) and B(58)) xor (A(122) and B(57)) xor (A(123) and B(56)) xor (A(124) and B(55)) xor (A(125) and B(54)) xor (A(126) and B(53)) xor (A(53) and B(127)) xor (A(54) and B(126)) xor (A(55) and B(125)) xor (A(56) and B(124)) xor (A(57) and B(123)) xor (A(58) and B(122)) xor (A(59) and B(121)) xor (A(60) and B(120)) xor (A(61) and B(119)) xor (A(62) and B(118)) xor (A(63) and B(117)) xor (A(64) and B(116)) xor (A(65) and B(115)) xor (A(66) and B(114)) xor (A(67) and B(113)) xor (A(68) and B(112)) xor (A(69) and B(111)) xor (A(70) and B(110)) xor (A(71) and B(109)) xor (A(72) and B(108)) xor (A(73) and B(107)) xor (A(74) and B(106)) xor (A(75) and B(105)) xor (A(76) and B(104)) xor (A(77) and B(103)) xor (A(78) and B(102)) xor (A(79) and B(101)) xor (A(80) and B(100)) xor (A(81) and B(99)) xor (A(82) and B(98)) xor (A(83) and B(97)) xor (A(84) and B(96)) xor (A(85) and B(95)) xor (A(86) and B(94)) xor (A(87) and B(93)) xor (A(88) and B(92)) xor (A(89) and B(91)) xor (A(90) and B(90)) xor (A(91) and B(89)) xor (A(92) and B(88)) xor (A(93) and B(87)) xor (A(94) and B(86)) xor (A(95) and B(85)) xor (A(96) and B(84)) xor (A(97) and B(83)) xor (A(98) and B(82)) xor (A(99) and B(81)) xor (A(100) and B(80)) xor (A(101) and B(79)) xor (A(102) and B(78)) xor (A(103) and B(77)) xor (A(104) and B(76)) xor (A(105) and B(75)) xor (A(106) and B(74)) xor (A(107) and B(73)) xor (A(108) and B(72)) xor (A(109) and B(71)) xor (A(110) and B(70)) xor (A(111) and B(69)) xor (A(112) and B(68)) xor (A(113) and B(67)) xor (A(114) and B(66)) xor (A(115) and B(65)) xor (A(116) and B(64)) xor (A(117) and B(63)) xor (A(118) and B(62)) xor (A(119) and B(61)) xor (A(120) and B(60)) xor (A(121) and B(59)) xor (A(122) and B(58)) xor (A(123) and B(57)) xor (A(124) and B(56)) xor (A(125) and B(55)) xor (A(126) and B(55));
    C(54)  <= (A(0) and B(54)) xor (A(1) and B(53)) xor (A(2) and B(52)) xor (A(3) and B(51)) xor (A(4) and B(50)) xor (A(5) and B(49)) xor (A(6) and B(48)) xor (A(7) and B(47)) xor (A(8) and B(46)) xor (A(9) and B(45)) xor (A(10) and B(44)) xor (A(11) and B(43)) xor (A(12) and B(42)) xor (A(13) and B(41)) xor (A(14) and B(40)) xor (A(15) and B(39)) xor (A(16) and B(38)) xor (A(17) and B(37)) xor (A(18) and B(36)) xor (A(19) and B(35)) xor (A(20) and B(34)) xor (A(21) and B(33)) xor (A(23) and B(32)) xor (A(23) and B(31)) xor (A(24) and B(30)) xor (A(25) and B(29)) xor (A(26) and B(28)) xor (A(27) and B(27)) xor (A(28) and B(26)) xor (A(29) and B(25)) xor (A(30) and B(24)) xor (A(31) and B(23)) xor (A(32) and B(23)) xor (A(33) and B(21)) xor (A(34) and B(20)) xor (A(35) and B(19)) xor (A(36) and B(18)) xor (A(37) and B(17)) xor (A(38) and B(16)) xor (A(39) and B(15)) xor (A(40) and B(14)) xor (A(41) and B(13)) xor (A(42) and B(12)) xor (A(43) and B(11)) xor (A(44) and B(10)) xor (A(45) and B(9)) xor (A(46) and B(8)) xor (A(47) and B(7)) xor (A(48) and B(6)) xor (A(49) and B(5)) xor (A(50) and B(4)) xor (A(51) and B(3)) xor (A(52) and B(2)) xor (A(53) and B(1)) xor (A(54) and B(0)) xor (A(47) and B(127)) xor (A(48) and B(126)) xor (A(49) and B(125)) xor (A(50) and B(124)) xor (A(51) and B(123)) xor (A(52) and B(122)) xor (A(53) and B(121)) xor (A(54) and B(120)) xor (A(55) and B(119)) xor (A(56) and B(118)) xor (A(57) and B(117)) xor (A(58) and B(116)) xor (A(59) and B(115)) xor (A(60) and B(114)) xor (A(61) and B(113)) xor (A(62) and B(112)) xor (A(63) and B(111)) xor (A(64) and B(110)) xor (A(65) and B(109)) xor (A(66) and B(108)) xor (A(67) and B(107)) xor (A(68) and B(106)) xor (A(69) and B(105)) xor (A(70) and B(104)) xor (A(71) and B(103)) xor (A(72) and B(102)) xor (A(73) and B(101)) xor (A(74) and B(100)) xor (A(75) and B(99)) xor (A(76) and B(98)) xor (A(77) and B(97)) xor (A(78) and B(96)) xor (A(79) and B(95)) xor (A(80) and B(94)) xor (A(81) and B(93)) xor (A(82) and B(92)) xor (A(83) and B(91)) xor (A(84) and B(90)) xor (A(85) and B(89)) xor (A(86) and B(88)) xor (A(87) and B(87)) xor (A(88) and B(86)) xor (A(89) and B(85)) xor (A(90) and B(84)) xor (A(91) and B(83)) xor (A(92) and B(82)) xor (A(93) and B(81)) xor (A(94) and B(80)) xor (A(95) and B(79)) xor (A(96) and B(78)) xor (A(97) and B(77)) xor (A(98) and B(76)) xor (A(99) and B(75)) xor (A(100) and B(74)) xor (A(101) and B(73)) xor (A(102) and B(72)) xor (A(103) and B(71)) xor (A(104) and B(70)) xor (A(105) and B(69)) xor (A(106) and B(68)) xor (A(107) and B(67)) xor (A(108) and B(66)) xor (A(109) and B(65)) xor (A(110) and B(64)) xor (A(111) and B(63)) xor (A(112) and B(62)) xor (A(113) and B(61)) xor (A(114) and B(60)) xor (A(115) and B(59)) xor (A(116) and B(58)) xor (A(117) and B(57)) xor (A(118) and B(56)) xor (A(119) and B(55)) xor (A(120) and B(54)) xor (A(121) and B(53)) xor (A(122) and B(52)) xor (A(123) and B(51)) xor (A(124) and B(50)) xor (A(125) and B(49)) xor (A(126) and B(48)) xor (A(52) and B(127)) xor (A(53) and B(126)) xor (A(54) and B(125)) xor (A(55) and B(124)) xor (A(56) and B(123)) xor (A(57) and B(122)) xor (A(58) and B(121)) xor (A(59) and B(120)) xor (A(60) and B(119)) xor (A(61) and B(118)) xor (A(62) and B(117)) xor (A(63) and B(116)) xor (A(64) and B(115)) xor (A(65) and B(114)) xor (A(66) and B(113)) xor (A(67) and B(112)) xor (A(68) and B(111)) xor (A(69) and B(110)) xor (A(70) and B(109)) xor (A(71) and B(108)) xor (A(72) and B(107)) xor (A(73) and B(106)) xor (A(74) and B(105)) xor (A(75) and B(104)) xor (A(76) and B(103)) xor (A(77) and B(102)) xor (A(78) and B(101)) xor (A(79) and B(100)) xor (A(80) and B(99)) xor (A(81) and B(98)) xor (A(82) and B(97)) xor (A(83) and B(96)) xor (A(84) and B(95)) xor (A(85) and B(94)) xor (A(86) and B(93)) xor (A(87) and B(92)) xor (A(88) and B(91)) xor (A(89) and B(90)) xor (A(90) and B(89)) xor (A(91) and B(88)) xor (A(92) and B(87)) xor (A(93) and B(86)) xor (A(94) and B(85)) xor (A(95) and B(84)) xor (A(96) and B(83)) xor (A(97) and B(82)) xor (A(98) and B(81)) xor (A(99) and B(80)) xor (A(100) and B(79)) xor (A(101) and B(78)) xor (A(102) and B(77)) xor (A(103) and B(76)) xor (A(104) and B(75)) xor (A(105) and B(74)) xor (A(106) and B(73)) xor (A(107) and B(72)) xor (A(108) and B(71)) xor (A(109) and B(70)) xor (A(110) and B(69)) xor (A(111) and B(68)) xor (A(112) and B(67)) xor (A(113) and B(66)) xor (A(114) and B(65)) xor (A(115) and B(64)) xor (A(116) and B(63)) xor (A(117) and B(62)) xor (A(118) and B(61)) xor (A(119) and B(60)) xor (A(120) and B(59)) xor (A(121) and B(58)) xor (A(122) and B(57)) xor (A(123) and B(56)) xor (A(124) and B(55)) xor (A(125) and B(54)) xor (A(126) and B(53)) xor (A(53) and B(127)) xor (A(54) and B(126)) xor (A(55) and B(125)) xor (A(56) and B(124)) xor (A(57) and B(123)) xor (A(58) and B(122)) xor (A(59) and B(121)) xor (A(60) and B(120)) xor (A(61) and B(119)) xor (A(62) and B(118)) xor (A(63) and B(117)) xor (A(64) and B(116)) xor (A(65) and B(115)) xor (A(66) and B(114)) xor (A(67) and B(113)) xor (A(68) and B(112)) xor (A(69) and B(111)) xor (A(70) and B(110)) xor (A(71) and B(109)) xor (A(72) and B(108)) xor (A(73) and B(107)) xor (A(74) and B(106)) xor (A(75) and B(105)) xor (A(76) and B(104)) xor (A(77) and B(103)) xor (A(78) and B(102)) xor (A(79) and B(101)) xor (A(80) and B(100)) xor (A(81) and B(99)) xor (A(82) and B(98)) xor (A(83) and B(97)) xor (A(84) and B(96)) xor (A(85) and B(95)) xor (A(86) and B(94)) xor (A(87) and B(93)) xor (A(88) and B(92)) xor (A(89) and B(91)) xor (A(90) and B(90)) xor (A(91) and B(89)) xor (A(92) and B(88)) xor (A(93) and B(87)) xor (A(94) and B(86)) xor (A(95) and B(85)) xor (A(96) and B(84)) xor (A(97) and B(83)) xor (A(98) and B(82)) xor (A(99) and B(81)) xor (A(100) and B(80)) xor (A(101) and B(79)) xor (A(102) and B(78)) xor (A(103) and B(77)) xor (A(104) and B(76)) xor (A(105) and B(75)) xor (A(106) and B(74)) xor (A(107) and B(73)) xor (A(108) and B(72)) xor (A(109) and B(71)) xor (A(110) and B(70)) xor (A(111) and B(69)) xor (A(112) and B(68)) xor (A(113) and B(67)) xor (A(114) and B(66)) xor (A(115) and B(65)) xor (A(116) and B(64)) xor (A(117) and B(63)) xor (A(118) and B(62)) xor (A(119) and B(61)) xor (A(120) and B(60)) xor (A(121) and B(59)) xor (A(122) and B(58)) xor (A(123) and B(57)) xor (A(124) and B(56)) xor (A(125) and B(55)) xor (A(126) and B(54)) xor (A(54) and B(127)) xor (A(55) and B(126)) xor (A(56) and B(125)) xor (A(57) and B(124)) xor (A(58) and B(123)) xor (A(59) and B(122)) xor (A(60) and B(121)) xor (A(61) and B(120)) xor (A(62) and B(119)) xor (A(63) and B(118)) xor (A(64) and B(117)) xor (A(65) and B(116)) xor (A(66) and B(115)) xor (A(67) and B(114)) xor (A(68) and B(113)) xor (A(69) and B(112)) xor (A(70) and B(111)) xor (A(71) and B(110)) xor (A(72) and B(109)) xor (A(73) and B(108)) xor (A(74) and B(107)) xor (A(75) and B(106)) xor (A(76) and B(105)) xor (A(77) and B(104)) xor (A(78) and B(103)) xor (A(79) and B(102)) xor (A(80) and B(101)) xor (A(81) and B(100)) xor (A(82) and B(99)) xor (A(83) and B(98)) xor (A(84) and B(97)) xor (A(85) and B(96)) xor (A(86) and B(95)) xor (A(87) and B(94)) xor (A(88) and B(93)) xor (A(89) and B(92)) xor (A(90) and B(91)) xor (A(91) and B(90)) xor (A(92) and B(89)) xor (A(93) and B(88)) xor (A(94) and B(87)) xor (A(95) and B(86)) xor (A(96) and B(85)) xor (A(97) and B(84)) xor (A(98) and B(83)) xor (A(99) and B(82)) xor (A(100) and B(81)) xor (A(101) and B(80)) xor (A(102) and B(79)) xor (A(103) and B(78)) xor (A(104) and B(77)) xor (A(105) and B(76)) xor (A(106) and B(75)) xor (A(107) and B(74)) xor (A(108) and B(73)) xor (A(109) and B(72)) xor (A(110) and B(71)) xor (A(111) and B(70)) xor (A(112) and B(69)) xor (A(113) and B(68)) xor (A(114) and B(67)) xor (A(115) and B(66)) xor (A(116) and B(65)) xor (A(117) and B(64)) xor (A(118) and B(63)) xor (A(119) and B(62)) xor (A(120) and B(61)) xor (A(121) and B(60)) xor (A(122) and B(59)) xor (A(123) and B(58)) xor (A(124) and B(57)) xor (A(125) and B(56)) xor (A(126) and B(56));
    C(55)  <= (A(0) and B(55)) xor (A(1) and B(54)) xor (A(2) and B(53)) xor (A(3) and B(52)) xor (A(4) and B(51)) xor (A(5) and B(50)) xor (A(6) and B(49)) xor (A(7) and B(48)) xor (A(8) and B(47)) xor (A(9) and B(46)) xor (A(10) and B(45)) xor (A(11) and B(44)) xor (A(12) and B(43)) xor (A(13) and B(42)) xor (A(14) and B(41)) xor (A(15) and B(40)) xor (A(16) and B(39)) xor (A(17) and B(38)) xor (A(18) and B(37)) xor (A(19) and B(36)) xor (A(20) and B(35)) xor (A(21) and B(34)) xor (A(23) and B(33)) xor (A(23) and B(32)) xor (A(24) and B(31)) xor (A(25) and B(30)) xor (A(26) and B(29)) xor (A(27) and B(28)) xor (A(28) and B(27)) xor (A(29) and B(26)) xor (A(30) and B(25)) xor (A(31) and B(24)) xor (A(32) and B(23)) xor (A(33) and B(23)) xor (A(34) and B(21)) xor (A(35) and B(20)) xor (A(36) and B(19)) xor (A(37) and B(18)) xor (A(38) and B(17)) xor (A(39) and B(16)) xor (A(40) and B(15)) xor (A(41) and B(14)) xor (A(42) and B(13)) xor (A(43) and B(12)) xor (A(44) and B(11)) xor (A(45) and B(10)) xor (A(46) and B(9)) xor (A(47) and B(8)) xor (A(48) and B(7)) xor (A(49) and B(6)) xor (A(50) and B(5)) xor (A(51) and B(4)) xor (A(52) and B(3)) xor (A(53) and B(2)) xor (A(54) and B(1)) xor (A(55) and B(0)) xor (A(48) and B(127)) xor (A(49) and B(126)) xor (A(50) and B(125)) xor (A(51) and B(124)) xor (A(52) and B(123)) xor (A(53) and B(122)) xor (A(54) and B(121)) xor (A(55) and B(120)) xor (A(56) and B(119)) xor (A(57) and B(118)) xor (A(58) and B(117)) xor (A(59) and B(116)) xor (A(60) and B(115)) xor (A(61) and B(114)) xor (A(62) and B(113)) xor (A(63) and B(112)) xor (A(64) and B(111)) xor (A(65) and B(110)) xor (A(66) and B(109)) xor (A(67) and B(108)) xor (A(68) and B(107)) xor (A(69) and B(106)) xor (A(70) and B(105)) xor (A(71) and B(104)) xor (A(72) and B(103)) xor (A(73) and B(102)) xor (A(74) and B(101)) xor (A(75) and B(100)) xor (A(76) and B(99)) xor (A(77) and B(98)) xor (A(78) and B(97)) xor (A(79) and B(96)) xor (A(80) and B(95)) xor (A(81) and B(94)) xor (A(82) and B(93)) xor (A(83) and B(92)) xor (A(84) and B(91)) xor (A(85) and B(90)) xor (A(86) and B(89)) xor (A(87) and B(88)) xor (A(88) and B(87)) xor (A(89) and B(86)) xor (A(90) and B(85)) xor (A(91) and B(84)) xor (A(92) and B(83)) xor (A(93) and B(82)) xor (A(94) and B(81)) xor (A(95) and B(80)) xor (A(96) and B(79)) xor (A(97) and B(78)) xor (A(98) and B(77)) xor (A(99) and B(76)) xor (A(100) and B(75)) xor (A(101) and B(74)) xor (A(102) and B(73)) xor (A(103) and B(72)) xor (A(104) and B(71)) xor (A(105) and B(70)) xor (A(106) and B(69)) xor (A(107) and B(68)) xor (A(108) and B(67)) xor (A(109) and B(66)) xor (A(110) and B(65)) xor (A(111) and B(64)) xor (A(112) and B(63)) xor (A(113) and B(62)) xor (A(114) and B(61)) xor (A(115) and B(60)) xor (A(116) and B(59)) xor (A(117) and B(58)) xor (A(118) and B(57)) xor (A(119) and B(56)) xor (A(120) and B(55)) xor (A(121) and B(54)) xor (A(122) and B(53)) xor (A(123) and B(52)) xor (A(124) and B(51)) xor (A(125) and B(50)) xor (A(126) and B(49)) xor (A(53) and B(127)) xor (A(54) and B(126)) xor (A(55) and B(125)) xor (A(56) and B(124)) xor (A(57) and B(123)) xor (A(58) and B(122)) xor (A(59) and B(121)) xor (A(60) and B(120)) xor (A(61) and B(119)) xor (A(62) and B(118)) xor (A(63) and B(117)) xor (A(64) and B(116)) xor (A(65) and B(115)) xor (A(66) and B(114)) xor (A(67) and B(113)) xor (A(68) and B(112)) xor (A(69) and B(111)) xor (A(70) and B(110)) xor (A(71) and B(109)) xor (A(72) and B(108)) xor (A(73) and B(107)) xor (A(74) and B(106)) xor (A(75) and B(105)) xor (A(76) and B(104)) xor (A(77) and B(103)) xor (A(78) and B(102)) xor (A(79) and B(101)) xor (A(80) and B(100)) xor (A(81) and B(99)) xor (A(82) and B(98)) xor (A(83) and B(97)) xor (A(84) and B(96)) xor (A(85) and B(95)) xor (A(86) and B(94)) xor (A(87) and B(93)) xor (A(88) and B(92)) xor (A(89) and B(91)) xor (A(90) and B(90)) xor (A(91) and B(89)) xor (A(92) and B(88)) xor (A(93) and B(87)) xor (A(94) and B(86)) xor (A(95) and B(85)) xor (A(96) and B(84)) xor (A(97) and B(83)) xor (A(98) and B(82)) xor (A(99) and B(81)) xor (A(100) and B(80)) xor (A(101) and B(79)) xor (A(102) and B(78)) xor (A(103) and B(77)) xor (A(104) and B(76)) xor (A(105) and B(75)) xor (A(106) and B(74)) xor (A(107) and B(73)) xor (A(108) and B(72)) xor (A(109) and B(71)) xor (A(110) and B(70)) xor (A(111) and B(69)) xor (A(112) and B(68)) xor (A(113) and B(67)) xor (A(114) and B(66)) xor (A(115) and B(65)) xor (A(116) and B(64)) xor (A(117) and B(63)) xor (A(118) and B(62)) xor (A(119) and B(61)) xor (A(120) and B(60)) xor (A(121) and B(59)) xor (A(122) and B(58)) xor (A(123) and B(57)) xor (A(124) and B(56)) xor (A(125) and B(55)) xor (A(126) and B(54)) xor (A(54) and B(127)) xor (A(55) and B(126)) xor (A(56) and B(125)) xor (A(57) and B(124)) xor (A(58) and B(123)) xor (A(59) and B(122)) xor (A(60) and B(121)) xor (A(61) and B(120)) xor (A(62) and B(119)) xor (A(63) and B(118)) xor (A(64) and B(117)) xor (A(65) and B(116)) xor (A(66) and B(115)) xor (A(67) and B(114)) xor (A(68) and B(113)) xor (A(69) and B(112)) xor (A(70) and B(111)) xor (A(71) and B(110)) xor (A(72) and B(109)) xor (A(73) and B(108)) xor (A(74) and B(107)) xor (A(75) and B(106)) xor (A(76) and B(105)) xor (A(77) and B(104)) xor (A(78) and B(103)) xor (A(79) and B(102)) xor (A(80) and B(101)) xor (A(81) and B(100)) xor (A(82) and B(99)) xor (A(83) and B(98)) xor (A(84) and B(97)) xor (A(85) and B(96)) xor (A(86) and B(95)) xor (A(87) and B(94)) xor (A(88) and B(93)) xor (A(89) and B(92)) xor (A(90) and B(91)) xor (A(91) and B(90)) xor (A(92) and B(89)) xor (A(93) and B(88)) xor (A(94) and B(87)) xor (A(95) and B(86)) xor (A(96) and B(85)) xor (A(97) and B(84)) xor (A(98) and B(83)) xor (A(99) and B(82)) xor (A(100) and B(81)) xor (A(101) and B(80)) xor (A(102) and B(79)) xor (A(103) and B(78)) xor (A(104) and B(77)) xor (A(105) and B(76)) xor (A(106) and B(75)) xor (A(107) and B(74)) xor (A(108) and B(73)) xor (A(109) and B(72)) xor (A(110) and B(71)) xor (A(111) and B(70)) xor (A(112) and B(69)) xor (A(113) and B(68)) xor (A(114) and B(67)) xor (A(115) and B(66)) xor (A(116) and B(65)) xor (A(117) and B(64)) xor (A(118) and B(63)) xor (A(119) and B(62)) xor (A(120) and B(61)) xor (A(121) and B(60)) xor (A(122) and B(59)) xor (A(123) and B(58)) xor (A(124) and B(57)) xor (A(125) and B(56)) xor (A(126) and B(55)) xor (A(55) and B(127)) xor (A(56) and B(126)) xor (A(57) and B(125)) xor (A(58) and B(124)) xor (A(59) and B(123)) xor (A(60) and B(122)) xor (A(61) and B(121)) xor (A(62) and B(120)) xor (A(63) and B(119)) xor (A(64) and B(118)) xor (A(65) and B(117)) xor (A(66) and B(116)) xor (A(67) and B(115)) xor (A(68) and B(114)) xor (A(69) and B(113)) xor (A(70) and B(112)) xor (A(71) and B(111)) xor (A(72) and B(110)) xor (A(73) and B(109)) xor (A(74) and B(108)) xor (A(75) and B(107)) xor (A(76) and B(106)) xor (A(77) and B(105)) xor (A(78) and B(104)) xor (A(79) and B(103)) xor (A(80) and B(102)) xor (A(81) and B(101)) xor (A(82) and B(100)) xor (A(83) and B(99)) xor (A(84) and B(98)) xor (A(85) and B(97)) xor (A(86) and B(96)) xor (A(87) and B(95)) xor (A(88) and B(94)) xor (A(89) and B(93)) xor (A(90) and B(92)) xor (A(91) and B(91)) xor (A(92) and B(90)) xor (A(93) and B(89)) xor (A(94) and B(88)) xor (A(95) and B(87)) xor (A(96) and B(86)) xor (A(97) and B(85)) xor (A(98) and B(84)) xor (A(99) and B(83)) xor (A(100) and B(82)) xor (A(101) and B(81)) xor (A(102) and B(80)) xor (A(103) and B(79)) xor (A(104) and B(78)) xor (A(105) and B(77)) xor (A(106) and B(76)) xor (A(107) and B(75)) xor (A(108) and B(74)) xor (A(109) and B(73)) xor (A(110) and B(72)) xor (A(111) and B(71)) xor (A(112) and B(70)) xor (A(113) and B(69)) xor (A(114) and B(68)) xor (A(115) and B(67)) xor (A(116) and B(66)) xor (A(117) and B(65)) xor (A(118) and B(64)) xor (A(119) and B(63)) xor (A(120) and B(62)) xor (A(121) and B(61)) xor (A(122) and B(60)) xor (A(123) and B(59)) xor (A(124) and B(58)) xor (A(125) and B(57)) xor (A(126) and B(57));
    C(56)  <= (A(0) and B(56)) xor (A(1) and B(55)) xor (A(2) and B(54)) xor (A(3) and B(53)) xor (A(4) and B(52)) xor (A(5) and B(51)) xor (A(6) and B(50)) xor (A(7) and B(49)) xor (A(8) and B(48)) xor (A(9) and B(47)) xor (A(10) and B(46)) xor (A(11) and B(45)) xor (A(12) and B(44)) xor (A(13) and B(43)) xor (A(14) and B(42)) xor (A(15) and B(41)) xor (A(16) and B(40)) xor (A(17) and B(39)) xor (A(18) and B(38)) xor (A(19) and B(37)) xor (A(20) and B(36)) xor (A(21) and B(35)) xor (A(23) and B(34)) xor (A(23) and B(33)) xor (A(24) and B(32)) xor (A(25) and B(31)) xor (A(26) and B(30)) xor (A(27) and B(29)) xor (A(28) and B(28)) xor (A(29) and B(27)) xor (A(30) and B(26)) xor (A(31) and B(25)) xor (A(32) and B(24)) xor (A(33) and B(23)) xor (A(34) and B(23)) xor (A(35) and B(21)) xor (A(36) and B(20)) xor (A(37) and B(19)) xor (A(38) and B(18)) xor (A(39) and B(17)) xor (A(40) and B(16)) xor (A(41) and B(15)) xor (A(42) and B(14)) xor (A(43) and B(13)) xor (A(44) and B(12)) xor (A(45) and B(11)) xor (A(46) and B(10)) xor (A(47) and B(9)) xor (A(48) and B(8)) xor (A(49) and B(7)) xor (A(50) and B(6)) xor (A(51) and B(5)) xor (A(52) and B(4)) xor (A(53) and B(3)) xor (A(54) and B(2)) xor (A(55) and B(1)) xor (A(56) and B(0)) xor (A(49) and B(127)) xor (A(50) and B(126)) xor (A(51) and B(125)) xor (A(52) and B(124)) xor (A(53) and B(123)) xor (A(54) and B(122)) xor (A(55) and B(121)) xor (A(56) and B(120)) xor (A(57) and B(119)) xor (A(58) and B(118)) xor (A(59) and B(117)) xor (A(60) and B(116)) xor (A(61) and B(115)) xor (A(62) and B(114)) xor (A(63) and B(113)) xor (A(64) and B(112)) xor (A(65) and B(111)) xor (A(66) and B(110)) xor (A(67) and B(109)) xor (A(68) and B(108)) xor (A(69) and B(107)) xor (A(70) and B(106)) xor (A(71) and B(105)) xor (A(72) and B(104)) xor (A(73) and B(103)) xor (A(74) and B(102)) xor (A(75) and B(101)) xor (A(76) and B(100)) xor (A(77) and B(99)) xor (A(78) and B(98)) xor (A(79) and B(97)) xor (A(80) and B(96)) xor (A(81) and B(95)) xor (A(82) and B(94)) xor (A(83) and B(93)) xor (A(84) and B(92)) xor (A(85) and B(91)) xor (A(86) and B(90)) xor (A(87) and B(89)) xor (A(88) and B(88)) xor (A(89) and B(87)) xor (A(90) and B(86)) xor (A(91) and B(85)) xor (A(92) and B(84)) xor (A(93) and B(83)) xor (A(94) and B(82)) xor (A(95) and B(81)) xor (A(96) and B(80)) xor (A(97) and B(79)) xor (A(98) and B(78)) xor (A(99) and B(77)) xor (A(100) and B(76)) xor (A(101) and B(75)) xor (A(102) and B(74)) xor (A(103) and B(73)) xor (A(104) and B(72)) xor (A(105) and B(71)) xor (A(106) and B(70)) xor (A(107) and B(69)) xor (A(108) and B(68)) xor (A(109) and B(67)) xor (A(110) and B(66)) xor (A(111) and B(65)) xor (A(112) and B(64)) xor (A(113) and B(63)) xor (A(114) and B(62)) xor (A(115) and B(61)) xor (A(116) and B(60)) xor (A(117) and B(59)) xor (A(118) and B(58)) xor (A(119) and B(57)) xor (A(120) and B(56)) xor (A(121) and B(55)) xor (A(122) and B(54)) xor (A(123) and B(53)) xor (A(124) and B(52)) xor (A(125) and B(51)) xor (A(126) and B(50)) xor (A(54) and B(127)) xor (A(55) and B(126)) xor (A(56) and B(125)) xor (A(57) and B(124)) xor (A(58) and B(123)) xor (A(59) and B(122)) xor (A(60) and B(121)) xor (A(61) and B(120)) xor (A(62) and B(119)) xor (A(63) and B(118)) xor (A(64) and B(117)) xor (A(65) and B(116)) xor (A(66) and B(115)) xor (A(67) and B(114)) xor (A(68) and B(113)) xor (A(69) and B(112)) xor (A(70) and B(111)) xor (A(71) and B(110)) xor (A(72) and B(109)) xor (A(73) and B(108)) xor (A(74) and B(107)) xor (A(75) and B(106)) xor (A(76) and B(105)) xor (A(77) and B(104)) xor (A(78) and B(103)) xor (A(79) and B(102)) xor (A(80) and B(101)) xor (A(81) and B(100)) xor (A(82) and B(99)) xor (A(83) and B(98)) xor (A(84) and B(97)) xor (A(85) and B(96)) xor (A(86) and B(95)) xor (A(87) and B(94)) xor (A(88) and B(93)) xor (A(89) and B(92)) xor (A(90) and B(91)) xor (A(91) and B(90)) xor (A(92) and B(89)) xor (A(93) and B(88)) xor (A(94) and B(87)) xor (A(95) and B(86)) xor (A(96) and B(85)) xor (A(97) and B(84)) xor (A(98) and B(83)) xor (A(99) and B(82)) xor (A(100) and B(81)) xor (A(101) and B(80)) xor (A(102) and B(79)) xor (A(103) and B(78)) xor (A(104) and B(77)) xor (A(105) and B(76)) xor (A(106) and B(75)) xor (A(107) and B(74)) xor (A(108) and B(73)) xor (A(109) and B(72)) xor (A(110) and B(71)) xor (A(111) and B(70)) xor (A(112) and B(69)) xor (A(113) and B(68)) xor (A(114) and B(67)) xor (A(115) and B(66)) xor (A(116) and B(65)) xor (A(117) and B(64)) xor (A(118) and B(63)) xor (A(119) and B(62)) xor (A(120) and B(61)) xor (A(121) and B(60)) xor (A(122) and B(59)) xor (A(123) and B(58)) xor (A(124) and B(57)) xor (A(125) and B(56)) xor (A(126) and B(55)) xor (A(55) and B(127)) xor (A(56) and B(126)) xor (A(57) and B(125)) xor (A(58) and B(124)) xor (A(59) and B(123)) xor (A(60) and B(122)) xor (A(61) and B(121)) xor (A(62) and B(120)) xor (A(63) and B(119)) xor (A(64) and B(118)) xor (A(65) and B(117)) xor (A(66) and B(116)) xor (A(67) and B(115)) xor (A(68) and B(114)) xor (A(69) and B(113)) xor (A(70) and B(112)) xor (A(71) and B(111)) xor (A(72) and B(110)) xor (A(73) and B(109)) xor (A(74) and B(108)) xor (A(75) and B(107)) xor (A(76) and B(106)) xor (A(77) and B(105)) xor (A(78) and B(104)) xor (A(79) and B(103)) xor (A(80) and B(102)) xor (A(81) and B(101)) xor (A(82) and B(100)) xor (A(83) and B(99)) xor (A(84) and B(98)) xor (A(85) and B(97)) xor (A(86) and B(96)) xor (A(87) and B(95)) xor (A(88) and B(94)) xor (A(89) and B(93)) xor (A(90) and B(92)) xor (A(91) and B(91)) xor (A(92) and B(90)) xor (A(93) and B(89)) xor (A(94) and B(88)) xor (A(95) and B(87)) xor (A(96) and B(86)) xor (A(97) and B(85)) xor (A(98) and B(84)) xor (A(99) and B(83)) xor (A(100) and B(82)) xor (A(101) and B(81)) xor (A(102) and B(80)) xor (A(103) and B(79)) xor (A(104) and B(78)) xor (A(105) and B(77)) xor (A(106) and B(76)) xor (A(107) and B(75)) xor (A(108) and B(74)) xor (A(109) and B(73)) xor (A(110) and B(72)) xor (A(111) and B(71)) xor (A(112) and B(70)) xor (A(113) and B(69)) xor (A(114) and B(68)) xor (A(115) and B(67)) xor (A(116) and B(66)) xor (A(117) and B(65)) xor (A(118) and B(64)) xor (A(119) and B(63)) xor (A(120) and B(62)) xor (A(121) and B(61)) xor (A(122) and B(60)) xor (A(123) and B(59)) xor (A(124) and B(58)) xor (A(125) and B(57)) xor (A(126) and B(56)) xor (A(56) and B(127)) xor (A(57) and B(126)) xor (A(58) and B(125)) xor (A(59) and B(124)) xor (A(60) and B(123)) xor (A(61) and B(122)) xor (A(62) and B(121)) xor (A(63) and B(120)) xor (A(64) and B(119)) xor (A(65) and B(118)) xor (A(66) and B(117)) xor (A(67) and B(116)) xor (A(68) and B(115)) xor (A(69) and B(114)) xor (A(70) and B(113)) xor (A(71) and B(112)) xor (A(72) and B(111)) xor (A(73) and B(110)) xor (A(74) and B(109)) xor (A(75) and B(108)) xor (A(76) and B(107)) xor (A(77) and B(106)) xor (A(78) and B(105)) xor (A(79) and B(104)) xor (A(80) and B(103)) xor (A(81) and B(102)) xor (A(82) and B(101)) xor (A(83) and B(100)) xor (A(84) and B(99)) xor (A(85) and B(98)) xor (A(86) and B(97)) xor (A(87) and B(96)) xor (A(88) and B(95)) xor (A(89) and B(94)) xor (A(90) and B(93)) xor (A(91) and B(92)) xor (A(92) and B(91)) xor (A(93) and B(90)) xor (A(94) and B(89)) xor (A(95) and B(88)) xor (A(96) and B(87)) xor (A(97) and B(86)) xor (A(98) and B(85)) xor (A(99) and B(84)) xor (A(100) and B(83)) xor (A(101) and B(82)) xor (A(102) and B(81)) xor (A(103) and B(80)) xor (A(104) and B(79)) xor (A(105) and B(78)) xor (A(106) and B(77)) xor (A(107) and B(76)) xor (A(108) and B(75)) xor (A(109) and B(74)) xor (A(110) and B(73)) xor (A(111) and B(72)) xor (A(112) and B(71)) xor (A(113) and B(70)) xor (A(114) and B(69)) xor (A(115) and B(68)) xor (A(116) and B(67)) xor (A(117) and B(66)) xor (A(118) and B(65)) xor (A(119) and B(64)) xor (A(120) and B(63)) xor (A(121) and B(62)) xor (A(122) and B(61)) xor (A(123) and B(60)) xor (A(124) and B(59)) xor (A(125) and B(58)) xor (A(126) and B(58));
    C(57)  <= (A(0) and B(57)) xor (A(1) and B(56)) xor (A(2) and B(55)) xor (A(3) and B(54)) xor (A(4) and B(53)) xor (A(5) and B(52)) xor (A(6) and B(51)) xor (A(7) and B(50)) xor (A(8) and B(49)) xor (A(9) and B(48)) xor (A(10) and B(47)) xor (A(11) and B(46)) xor (A(12) and B(45)) xor (A(13) and B(44)) xor (A(14) and B(43)) xor (A(15) and B(42)) xor (A(16) and B(41)) xor (A(17) and B(40)) xor (A(18) and B(39)) xor (A(19) and B(38)) xor (A(20) and B(37)) xor (A(21) and B(36)) xor (A(23) and B(35)) xor (A(23) and B(34)) xor (A(24) and B(33)) xor (A(25) and B(32)) xor (A(26) and B(31)) xor (A(27) and B(30)) xor (A(28) and B(29)) xor (A(29) and B(28)) xor (A(30) and B(27)) xor (A(31) and B(26)) xor (A(32) and B(25)) xor (A(33) and B(24)) xor (A(34) and B(23)) xor (A(35) and B(23)) xor (A(36) and B(21)) xor (A(37) and B(20)) xor (A(38) and B(19)) xor (A(39) and B(18)) xor (A(40) and B(17)) xor (A(41) and B(16)) xor (A(42) and B(15)) xor (A(43) and B(14)) xor (A(44) and B(13)) xor (A(45) and B(12)) xor (A(46) and B(11)) xor (A(47) and B(10)) xor (A(48) and B(9)) xor (A(49) and B(8)) xor (A(50) and B(7)) xor (A(51) and B(6)) xor (A(52) and B(5)) xor (A(53) and B(4)) xor (A(54) and B(3)) xor (A(55) and B(2)) xor (A(56) and B(1)) xor (A(57) and B(0)) xor (A(50) and B(127)) xor (A(51) and B(126)) xor (A(52) and B(125)) xor (A(53) and B(124)) xor (A(54) and B(123)) xor (A(55) and B(122)) xor (A(56) and B(121)) xor (A(57) and B(120)) xor (A(58) and B(119)) xor (A(59) and B(118)) xor (A(60) and B(117)) xor (A(61) and B(116)) xor (A(62) and B(115)) xor (A(63) and B(114)) xor (A(64) and B(113)) xor (A(65) and B(112)) xor (A(66) and B(111)) xor (A(67) and B(110)) xor (A(68) and B(109)) xor (A(69) and B(108)) xor (A(70) and B(107)) xor (A(71) and B(106)) xor (A(72) and B(105)) xor (A(73) and B(104)) xor (A(74) and B(103)) xor (A(75) and B(102)) xor (A(76) and B(101)) xor (A(77) and B(100)) xor (A(78) and B(99)) xor (A(79) and B(98)) xor (A(80) and B(97)) xor (A(81) and B(96)) xor (A(82) and B(95)) xor (A(83) and B(94)) xor (A(84) and B(93)) xor (A(85) and B(92)) xor (A(86) and B(91)) xor (A(87) and B(90)) xor (A(88) and B(89)) xor (A(89) and B(88)) xor (A(90) and B(87)) xor (A(91) and B(86)) xor (A(92) and B(85)) xor (A(93) and B(84)) xor (A(94) and B(83)) xor (A(95) and B(82)) xor (A(96) and B(81)) xor (A(97) and B(80)) xor (A(98) and B(79)) xor (A(99) and B(78)) xor (A(100) and B(77)) xor (A(101) and B(76)) xor (A(102) and B(75)) xor (A(103) and B(74)) xor (A(104) and B(73)) xor (A(105) and B(72)) xor (A(106) and B(71)) xor (A(107) and B(70)) xor (A(108) and B(69)) xor (A(109) and B(68)) xor (A(110) and B(67)) xor (A(111) and B(66)) xor (A(112) and B(65)) xor (A(113) and B(64)) xor (A(114) and B(63)) xor (A(115) and B(62)) xor (A(116) and B(61)) xor (A(117) and B(60)) xor (A(118) and B(59)) xor (A(119) and B(58)) xor (A(120) and B(57)) xor (A(121) and B(56)) xor (A(122) and B(55)) xor (A(123) and B(54)) xor (A(124) and B(53)) xor (A(125) and B(52)) xor (A(126) and B(51)) xor (A(55) and B(127)) xor (A(56) and B(126)) xor (A(57) and B(125)) xor (A(58) and B(124)) xor (A(59) and B(123)) xor (A(60) and B(122)) xor (A(61) and B(121)) xor (A(62) and B(120)) xor (A(63) and B(119)) xor (A(64) and B(118)) xor (A(65) and B(117)) xor (A(66) and B(116)) xor (A(67) and B(115)) xor (A(68) and B(114)) xor (A(69) and B(113)) xor (A(70) and B(112)) xor (A(71) and B(111)) xor (A(72) and B(110)) xor (A(73) and B(109)) xor (A(74) and B(108)) xor (A(75) and B(107)) xor (A(76) and B(106)) xor (A(77) and B(105)) xor (A(78) and B(104)) xor (A(79) and B(103)) xor (A(80) and B(102)) xor (A(81) and B(101)) xor (A(82) and B(100)) xor (A(83) and B(99)) xor (A(84) and B(98)) xor (A(85) and B(97)) xor (A(86) and B(96)) xor (A(87) and B(95)) xor (A(88) and B(94)) xor (A(89) and B(93)) xor (A(90) and B(92)) xor (A(91) and B(91)) xor (A(92) and B(90)) xor (A(93) and B(89)) xor (A(94) and B(88)) xor (A(95) and B(87)) xor (A(96) and B(86)) xor (A(97) and B(85)) xor (A(98) and B(84)) xor (A(99) and B(83)) xor (A(100) and B(82)) xor (A(101) and B(81)) xor (A(102) and B(80)) xor (A(103) and B(79)) xor (A(104) and B(78)) xor (A(105) and B(77)) xor (A(106) and B(76)) xor (A(107) and B(75)) xor (A(108) and B(74)) xor (A(109) and B(73)) xor (A(110) and B(72)) xor (A(111) and B(71)) xor (A(112) and B(70)) xor (A(113) and B(69)) xor (A(114) and B(68)) xor (A(115) and B(67)) xor (A(116) and B(66)) xor (A(117) and B(65)) xor (A(118) and B(64)) xor (A(119) and B(63)) xor (A(120) and B(62)) xor (A(121) and B(61)) xor (A(122) and B(60)) xor (A(123) and B(59)) xor (A(124) and B(58)) xor (A(125) and B(57)) xor (A(126) and B(56)) xor (A(56) and B(127)) xor (A(57) and B(126)) xor (A(58) and B(125)) xor (A(59) and B(124)) xor (A(60) and B(123)) xor (A(61) and B(122)) xor (A(62) and B(121)) xor (A(63) and B(120)) xor (A(64) and B(119)) xor (A(65) and B(118)) xor (A(66) and B(117)) xor (A(67) and B(116)) xor (A(68) and B(115)) xor (A(69) and B(114)) xor (A(70) and B(113)) xor (A(71) and B(112)) xor (A(72) and B(111)) xor (A(73) and B(110)) xor (A(74) and B(109)) xor (A(75) and B(108)) xor (A(76) and B(107)) xor (A(77) and B(106)) xor (A(78) and B(105)) xor (A(79) and B(104)) xor (A(80) and B(103)) xor (A(81) and B(102)) xor (A(82) and B(101)) xor (A(83) and B(100)) xor (A(84) and B(99)) xor (A(85) and B(98)) xor (A(86) and B(97)) xor (A(87) and B(96)) xor (A(88) and B(95)) xor (A(89) and B(94)) xor (A(90) and B(93)) xor (A(91) and B(92)) xor (A(92) and B(91)) xor (A(93) and B(90)) xor (A(94) and B(89)) xor (A(95) and B(88)) xor (A(96) and B(87)) xor (A(97) and B(86)) xor (A(98) and B(85)) xor (A(99) and B(84)) xor (A(100) and B(83)) xor (A(101) and B(82)) xor (A(102) and B(81)) xor (A(103) and B(80)) xor (A(104) and B(79)) xor (A(105) and B(78)) xor (A(106) and B(77)) xor (A(107) and B(76)) xor (A(108) and B(75)) xor (A(109) and B(74)) xor (A(110) and B(73)) xor (A(111) and B(72)) xor (A(112) and B(71)) xor (A(113) and B(70)) xor (A(114) and B(69)) xor (A(115) and B(68)) xor (A(116) and B(67)) xor (A(117) and B(66)) xor (A(118) and B(65)) xor (A(119) and B(64)) xor (A(120) and B(63)) xor (A(121) and B(62)) xor (A(122) and B(61)) xor (A(123) and B(60)) xor (A(124) and B(59)) xor (A(125) and B(58)) xor (A(126) and B(57)) xor (A(57) and B(127)) xor (A(58) and B(126)) xor (A(59) and B(125)) xor (A(60) and B(124)) xor (A(61) and B(123)) xor (A(62) and B(122)) xor (A(63) and B(121)) xor (A(64) and B(120)) xor (A(65) and B(119)) xor (A(66) and B(118)) xor (A(67) and B(117)) xor (A(68) and B(116)) xor (A(69) and B(115)) xor (A(70) and B(114)) xor (A(71) and B(113)) xor (A(72) and B(112)) xor (A(73) and B(111)) xor (A(74) and B(110)) xor (A(75) and B(109)) xor (A(76) and B(108)) xor (A(77) and B(107)) xor (A(78) and B(106)) xor (A(79) and B(105)) xor (A(80) and B(104)) xor (A(81) and B(103)) xor (A(82) and B(102)) xor (A(83) and B(101)) xor (A(84) and B(100)) xor (A(85) and B(99)) xor (A(86) and B(98)) xor (A(87) and B(97)) xor (A(88) and B(96)) xor (A(89) and B(95)) xor (A(90) and B(94)) xor (A(91) and B(93)) xor (A(92) and B(92)) xor (A(93) and B(91)) xor (A(94) and B(90)) xor (A(95) and B(89)) xor (A(96) and B(88)) xor (A(97) and B(87)) xor (A(98) and B(86)) xor (A(99) and B(85)) xor (A(100) and B(84)) xor (A(101) and B(83)) xor (A(102) and B(82)) xor (A(103) and B(81)) xor (A(104) and B(80)) xor (A(105) and B(79)) xor (A(106) and B(78)) xor (A(107) and B(77)) xor (A(108) and B(76)) xor (A(109) and B(75)) xor (A(110) and B(74)) xor (A(111) and B(73)) xor (A(112) and B(72)) xor (A(113) and B(71)) xor (A(114) and B(70)) xor (A(115) and B(69)) xor (A(116) and B(68)) xor (A(117) and B(67)) xor (A(118) and B(66)) xor (A(119) and B(65)) xor (A(120) and B(64)) xor (A(121) and B(63)) xor (A(122) and B(62)) xor (A(123) and B(61)) xor (A(124) and B(60)) xor (A(125) and B(59)) xor (A(126) and B(59));
    C(58)  <= (A(0) and B(58)) xor (A(1) and B(57)) xor (A(2) and B(56)) xor (A(3) and B(55)) xor (A(4) and B(54)) xor (A(5) and B(53)) xor (A(6) and B(52)) xor (A(7) and B(51)) xor (A(8) and B(50)) xor (A(9) and B(49)) xor (A(10) and B(48)) xor (A(11) and B(47)) xor (A(12) and B(46)) xor (A(13) and B(45)) xor (A(14) and B(44)) xor (A(15) and B(43)) xor (A(16) and B(42)) xor (A(17) and B(41)) xor (A(18) and B(40)) xor (A(19) and B(39)) xor (A(20) and B(38)) xor (A(21) and B(37)) xor (A(23) and B(36)) xor (A(23) and B(35)) xor (A(24) and B(34)) xor (A(25) and B(33)) xor (A(26) and B(32)) xor (A(27) and B(31)) xor (A(28) and B(30)) xor (A(29) and B(29)) xor (A(30) and B(28)) xor (A(31) and B(27)) xor (A(32) and B(26)) xor (A(33) and B(25)) xor (A(34) and B(24)) xor (A(35) and B(23)) xor (A(36) and B(23)) xor (A(37) and B(21)) xor (A(38) and B(20)) xor (A(39) and B(19)) xor (A(40) and B(18)) xor (A(41) and B(17)) xor (A(42) and B(16)) xor (A(43) and B(15)) xor (A(44) and B(14)) xor (A(45) and B(13)) xor (A(46) and B(12)) xor (A(47) and B(11)) xor (A(48) and B(10)) xor (A(49) and B(9)) xor (A(50) and B(8)) xor (A(51) and B(7)) xor (A(52) and B(6)) xor (A(53) and B(5)) xor (A(54) and B(4)) xor (A(55) and B(3)) xor (A(56) and B(2)) xor (A(57) and B(1)) xor (A(58) and B(0)) xor (A(51) and B(127)) xor (A(52) and B(126)) xor (A(53) and B(125)) xor (A(54) and B(124)) xor (A(55) and B(123)) xor (A(56) and B(122)) xor (A(57) and B(121)) xor (A(58) and B(120)) xor (A(59) and B(119)) xor (A(60) and B(118)) xor (A(61) and B(117)) xor (A(62) and B(116)) xor (A(63) and B(115)) xor (A(64) and B(114)) xor (A(65) and B(113)) xor (A(66) and B(112)) xor (A(67) and B(111)) xor (A(68) and B(110)) xor (A(69) and B(109)) xor (A(70) and B(108)) xor (A(71) and B(107)) xor (A(72) and B(106)) xor (A(73) and B(105)) xor (A(74) and B(104)) xor (A(75) and B(103)) xor (A(76) and B(102)) xor (A(77) and B(101)) xor (A(78) and B(100)) xor (A(79) and B(99)) xor (A(80) and B(98)) xor (A(81) and B(97)) xor (A(82) and B(96)) xor (A(83) and B(95)) xor (A(84) and B(94)) xor (A(85) and B(93)) xor (A(86) and B(92)) xor (A(87) and B(91)) xor (A(88) and B(90)) xor (A(89) and B(89)) xor (A(90) and B(88)) xor (A(91) and B(87)) xor (A(92) and B(86)) xor (A(93) and B(85)) xor (A(94) and B(84)) xor (A(95) and B(83)) xor (A(96) and B(82)) xor (A(97) and B(81)) xor (A(98) and B(80)) xor (A(99) and B(79)) xor (A(100) and B(78)) xor (A(101) and B(77)) xor (A(102) and B(76)) xor (A(103) and B(75)) xor (A(104) and B(74)) xor (A(105) and B(73)) xor (A(106) and B(72)) xor (A(107) and B(71)) xor (A(108) and B(70)) xor (A(109) and B(69)) xor (A(110) and B(68)) xor (A(111) and B(67)) xor (A(112) and B(66)) xor (A(113) and B(65)) xor (A(114) and B(64)) xor (A(115) and B(63)) xor (A(116) and B(62)) xor (A(117) and B(61)) xor (A(118) and B(60)) xor (A(119) and B(59)) xor (A(120) and B(58)) xor (A(121) and B(57)) xor (A(122) and B(56)) xor (A(123) and B(55)) xor (A(124) and B(54)) xor (A(125) and B(53)) xor (A(126) and B(52)) xor (A(56) and B(127)) xor (A(57) and B(126)) xor (A(58) and B(125)) xor (A(59) and B(124)) xor (A(60) and B(123)) xor (A(61) and B(122)) xor (A(62) and B(121)) xor (A(63) and B(120)) xor (A(64) and B(119)) xor (A(65) and B(118)) xor (A(66) and B(117)) xor (A(67) and B(116)) xor (A(68) and B(115)) xor (A(69) and B(114)) xor (A(70) and B(113)) xor (A(71) and B(112)) xor (A(72) and B(111)) xor (A(73) and B(110)) xor (A(74) and B(109)) xor (A(75) and B(108)) xor (A(76) and B(107)) xor (A(77) and B(106)) xor (A(78) and B(105)) xor (A(79) and B(104)) xor (A(80) and B(103)) xor (A(81) and B(102)) xor (A(82) and B(101)) xor (A(83) and B(100)) xor (A(84) and B(99)) xor (A(85) and B(98)) xor (A(86) and B(97)) xor (A(87) and B(96)) xor (A(88) and B(95)) xor (A(89) and B(94)) xor (A(90) and B(93)) xor (A(91) and B(92)) xor (A(92) and B(91)) xor (A(93) and B(90)) xor (A(94) and B(89)) xor (A(95) and B(88)) xor (A(96) and B(87)) xor (A(97) and B(86)) xor (A(98) and B(85)) xor (A(99) and B(84)) xor (A(100) and B(83)) xor (A(101) and B(82)) xor (A(102) and B(81)) xor (A(103) and B(80)) xor (A(104) and B(79)) xor (A(105) and B(78)) xor (A(106) and B(77)) xor (A(107) and B(76)) xor (A(108) and B(75)) xor (A(109) and B(74)) xor (A(110) and B(73)) xor (A(111) and B(72)) xor (A(112) and B(71)) xor (A(113) and B(70)) xor (A(114) and B(69)) xor (A(115) and B(68)) xor (A(116) and B(67)) xor (A(117) and B(66)) xor (A(118) and B(65)) xor (A(119) and B(64)) xor (A(120) and B(63)) xor (A(121) and B(62)) xor (A(122) and B(61)) xor (A(123) and B(60)) xor (A(124) and B(59)) xor (A(125) and B(58)) xor (A(126) and B(57)) xor (A(57) and B(127)) xor (A(58) and B(126)) xor (A(59) and B(125)) xor (A(60) and B(124)) xor (A(61) and B(123)) xor (A(62) and B(122)) xor (A(63) and B(121)) xor (A(64) and B(120)) xor (A(65) and B(119)) xor (A(66) and B(118)) xor (A(67) and B(117)) xor (A(68) and B(116)) xor (A(69) and B(115)) xor (A(70) and B(114)) xor (A(71) and B(113)) xor (A(72) and B(112)) xor (A(73) and B(111)) xor (A(74) and B(110)) xor (A(75) and B(109)) xor (A(76) and B(108)) xor (A(77) and B(107)) xor (A(78) and B(106)) xor (A(79) and B(105)) xor (A(80) and B(104)) xor (A(81) and B(103)) xor (A(82) and B(102)) xor (A(83) and B(101)) xor (A(84) and B(100)) xor (A(85) and B(99)) xor (A(86) and B(98)) xor (A(87) and B(97)) xor (A(88) and B(96)) xor (A(89) and B(95)) xor (A(90) and B(94)) xor (A(91) and B(93)) xor (A(92) and B(92)) xor (A(93) and B(91)) xor (A(94) and B(90)) xor (A(95) and B(89)) xor (A(96) and B(88)) xor (A(97) and B(87)) xor (A(98) and B(86)) xor (A(99) and B(85)) xor (A(100) and B(84)) xor (A(101) and B(83)) xor (A(102) and B(82)) xor (A(103) and B(81)) xor (A(104) and B(80)) xor (A(105) and B(79)) xor (A(106) and B(78)) xor (A(107) and B(77)) xor (A(108) and B(76)) xor (A(109) and B(75)) xor (A(110) and B(74)) xor (A(111) and B(73)) xor (A(112) and B(72)) xor (A(113) and B(71)) xor (A(114) and B(70)) xor (A(115) and B(69)) xor (A(116) and B(68)) xor (A(117) and B(67)) xor (A(118) and B(66)) xor (A(119) and B(65)) xor (A(120) and B(64)) xor (A(121) and B(63)) xor (A(122) and B(62)) xor (A(123) and B(61)) xor (A(124) and B(60)) xor (A(125) and B(59)) xor (A(126) and B(58)) xor (A(58) and B(127)) xor (A(59) and B(126)) xor (A(60) and B(125)) xor (A(61) and B(124)) xor (A(62) and B(123)) xor (A(63) and B(122)) xor (A(64) and B(121)) xor (A(65) and B(120)) xor (A(66) and B(119)) xor (A(67) and B(118)) xor (A(68) and B(117)) xor (A(69) and B(116)) xor (A(70) and B(115)) xor (A(71) and B(114)) xor (A(72) and B(113)) xor (A(73) and B(112)) xor (A(74) and B(111)) xor (A(75) and B(110)) xor (A(76) and B(109)) xor (A(77) and B(108)) xor (A(78) and B(107)) xor (A(79) and B(106)) xor (A(80) and B(105)) xor (A(81) and B(104)) xor (A(82) and B(103)) xor (A(83) and B(102)) xor (A(84) and B(101)) xor (A(85) and B(100)) xor (A(86) and B(99)) xor (A(87) and B(98)) xor (A(88) and B(97)) xor (A(89) and B(96)) xor (A(90) and B(95)) xor (A(91) and B(94)) xor (A(92) and B(93)) xor (A(93) and B(92)) xor (A(94) and B(91)) xor (A(95) and B(90)) xor (A(96) and B(89)) xor (A(97) and B(88)) xor (A(98) and B(87)) xor (A(99) and B(86)) xor (A(100) and B(85)) xor (A(101) and B(84)) xor (A(102) and B(83)) xor (A(103) and B(82)) xor (A(104) and B(81)) xor (A(105) and B(80)) xor (A(106) and B(79)) xor (A(107) and B(78)) xor (A(108) and B(77)) xor (A(109) and B(76)) xor (A(110) and B(75)) xor (A(111) and B(74)) xor (A(112) and B(73)) xor (A(113) and B(72)) xor (A(114) and B(71)) xor (A(115) and B(70)) xor (A(116) and B(69)) xor (A(117) and B(68)) xor (A(118) and B(67)) xor (A(119) and B(66)) xor (A(120) and B(65)) xor (A(121) and B(64)) xor (A(122) and B(63)) xor (A(123) and B(62)) xor (A(124) and B(61)) xor (A(125) and B(60)) xor (A(126) and B(60));
    C(59)  <= (A(0) and B(59)) xor (A(1) and B(58)) xor (A(2) and B(57)) xor (A(3) and B(56)) xor (A(4) and B(55)) xor (A(5) and B(54)) xor (A(6) and B(53)) xor (A(7) and B(52)) xor (A(8) and B(51)) xor (A(9) and B(50)) xor (A(10) and B(49)) xor (A(11) and B(48)) xor (A(12) and B(47)) xor (A(13) and B(46)) xor (A(14) and B(45)) xor (A(15) and B(44)) xor (A(16) and B(43)) xor (A(17) and B(42)) xor (A(18) and B(41)) xor (A(19) and B(40)) xor (A(20) and B(39)) xor (A(21) and B(38)) xor (A(23) and B(37)) xor (A(23) and B(36)) xor (A(24) and B(35)) xor (A(25) and B(34)) xor (A(26) and B(33)) xor (A(27) and B(32)) xor (A(28) and B(31)) xor (A(29) and B(30)) xor (A(30) and B(29)) xor (A(31) and B(28)) xor (A(32) and B(27)) xor (A(33) and B(26)) xor (A(34) and B(25)) xor (A(35) and B(24)) xor (A(36) and B(23)) xor (A(37) and B(23)) xor (A(38) and B(21)) xor (A(39) and B(20)) xor (A(40) and B(19)) xor (A(41) and B(18)) xor (A(42) and B(17)) xor (A(43) and B(16)) xor (A(44) and B(15)) xor (A(45) and B(14)) xor (A(46) and B(13)) xor (A(47) and B(12)) xor (A(48) and B(11)) xor (A(49) and B(10)) xor (A(50) and B(9)) xor (A(51) and B(8)) xor (A(52) and B(7)) xor (A(53) and B(6)) xor (A(54) and B(5)) xor (A(55) and B(4)) xor (A(56) and B(3)) xor (A(57) and B(2)) xor (A(58) and B(1)) xor (A(59) and B(0)) xor (A(52) and B(127)) xor (A(53) and B(126)) xor (A(54) and B(125)) xor (A(55) and B(124)) xor (A(56) and B(123)) xor (A(57) and B(122)) xor (A(58) and B(121)) xor (A(59) and B(120)) xor (A(60) and B(119)) xor (A(61) and B(118)) xor (A(62) and B(117)) xor (A(63) and B(116)) xor (A(64) and B(115)) xor (A(65) and B(114)) xor (A(66) and B(113)) xor (A(67) and B(112)) xor (A(68) and B(111)) xor (A(69) and B(110)) xor (A(70) and B(109)) xor (A(71) and B(108)) xor (A(72) and B(107)) xor (A(73) and B(106)) xor (A(74) and B(105)) xor (A(75) and B(104)) xor (A(76) and B(103)) xor (A(77) and B(102)) xor (A(78) and B(101)) xor (A(79) and B(100)) xor (A(80) and B(99)) xor (A(81) and B(98)) xor (A(82) and B(97)) xor (A(83) and B(96)) xor (A(84) and B(95)) xor (A(85) and B(94)) xor (A(86) and B(93)) xor (A(87) and B(92)) xor (A(88) and B(91)) xor (A(89) and B(90)) xor (A(90) and B(89)) xor (A(91) and B(88)) xor (A(92) and B(87)) xor (A(93) and B(86)) xor (A(94) and B(85)) xor (A(95) and B(84)) xor (A(96) and B(83)) xor (A(97) and B(82)) xor (A(98) and B(81)) xor (A(99) and B(80)) xor (A(100) and B(79)) xor (A(101) and B(78)) xor (A(102) and B(77)) xor (A(103) and B(76)) xor (A(104) and B(75)) xor (A(105) and B(74)) xor (A(106) and B(73)) xor (A(107) and B(72)) xor (A(108) and B(71)) xor (A(109) and B(70)) xor (A(110) and B(69)) xor (A(111) and B(68)) xor (A(112) and B(67)) xor (A(113) and B(66)) xor (A(114) and B(65)) xor (A(115) and B(64)) xor (A(116) and B(63)) xor (A(117) and B(62)) xor (A(118) and B(61)) xor (A(119) and B(60)) xor (A(120) and B(59)) xor (A(121) and B(58)) xor (A(122) and B(57)) xor (A(123) and B(56)) xor (A(124) and B(55)) xor (A(125) and B(54)) xor (A(126) and B(53)) xor (A(57) and B(127)) xor (A(58) and B(126)) xor (A(59) and B(125)) xor (A(60) and B(124)) xor (A(61) and B(123)) xor (A(62) and B(122)) xor (A(63) and B(121)) xor (A(64) and B(120)) xor (A(65) and B(119)) xor (A(66) and B(118)) xor (A(67) and B(117)) xor (A(68) and B(116)) xor (A(69) and B(115)) xor (A(70) and B(114)) xor (A(71) and B(113)) xor (A(72) and B(112)) xor (A(73) and B(111)) xor (A(74) and B(110)) xor (A(75) and B(109)) xor (A(76) and B(108)) xor (A(77) and B(107)) xor (A(78) and B(106)) xor (A(79) and B(105)) xor (A(80) and B(104)) xor (A(81) and B(103)) xor (A(82) and B(102)) xor (A(83) and B(101)) xor (A(84) and B(100)) xor (A(85) and B(99)) xor (A(86) and B(98)) xor (A(87) and B(97)) xor (A(88) and B(96)) xor (A(89) and B(95)) xor (A(90) and B(94)) xor (A(91) and B(93)) xor (A(92) and B(92)) xor (A(93) and B(91)) xor (A(94) and B(90)) xor (A(95) and B(89)) xor (A(96) and B(88)) xor (A(97) and B(87)) xor (A(98) and B(86)) xor (A(99) and B(85)) xor (A(100) and B(84)) xor (A(101) and B(83)) xor (A(102) and B(82)) xor (A(103) and B(81)) xor (A(104) and B(80)) xor (A(105) and B(79)) xor (A(106) and B(78)) xor (A(107) and B(77)) xor (A(108) and B(76)) xor (A(109) and B(75)) xor (A(110) and B(74)) xor (A(111) and B(73)) xor (A(112) and B(72)) xor (A(113) and B(71)) xor (A(114) and B(70)) xor (A(115) and B(69)) xor (A(116) and B(68)) xor (A(117) and B(67)) xor (A(118) and B(66)) xor (A(119) and B(65)) xor (A(120) and B(64)) xor (A(121) and B(63)) xor (A(122) and B(62)) xor (A(123) and B(61)) xor (A(124) and B(60)) xor (A(125) and B(59)) xor (A(126) and B(58)) xor (A(58) and B(127)) xor (A(59) and B(126)) xor (A(60) and B(125)) xor (A(61) and B(124)) xor (A(62) and B(123)) xor (A(63) and B(122)) xor (A(64) and B(121)) xor (A(65) and B(120)) xor (A(66) and B(119)) xor (A(67) and B(118)) xor (A(68) and B(117)) xor (A(69) and B(116)) xor (A(70) and B(115)) xor (A(71) and B(114)) xor (A(72) and B(113)) xor (A(73) and B(112)) xor (A(74) and B(111)) xor (A(75) and B(110)) xor (A(76) and B(109)) xor (A(77) and B(108)) xor (A(78) and B(107)) xor (A(79) and B(106)) xor (A(80) and B(105)) xor (A(81) and B(104)) xor (A(82) and B(103)) xor (A(83) and B(102)) xor (A(84) and B(101)) xor (A(85) and B(100)) xor (A(86) and B(99)) xor (A(87) and B(98)) xor (A(88) and B(97)) xor (A(89) and B(96)) xor (A(90) and B(95)) xor (A(91) and B(94)) xor (A(92) and B(93)) xor (A(93) and B(92)) xor (A(94) and B(91)) xor (A(95) and B(90)) xor (A(96) and B(89)) xor (A(97) and B(88)) xor (A(98) and B(87)) xor (A(99) and B(86)) xor (A(100) and B(85)) xor (A(101) and B(84)) xor (A(102) and B(83)) xor (A(103) and B(82)) xor (A(104) and B(81)) xor (A(105) and B(80)) xor (A(106) and B(79)) xor (A(107) and B(78)) xor (A(108) and B(77)) xor (A(109) and B(76)) xor (A(110) and B(75)) xor (A(111) and B(74)) xor (A(112) and B(73)) xor (A(113) and B(72)) xor (A(114) and B(71)) xor (A(115) and B(70)) xor (A(116) and B(69)) xor (A(117) and B(68)) xor (A(118) and B(67)) xor (A(119) and B(66)) xor (A(120) and B(65)) xor (A(121) and B(64)) xor (A(122) and B(63)) xor (A(123) and B(62)) xor (A(124) and B(61)) xor (A(125) and B(60)) xor (A(126) and B(59)) xor (A(59) and B(127)) xor (A(60) and B(126)) xor (A(61) and B(125)) xor (A(62) and B(124)) xor (A(63) and B(123)) xor (A(64) and B(122)) xor (A(65) and B(121)) xor (A(66) and B(120)) xor (A(67) and B(119)) xor (A(68) and B(118)) xor (A(69) and B(117)) xor (A(70) and B(116)) xor (A(71) and B(115)) xor (A(72) and B(114)) xor (A(73) and B(113)) xor (A(74) and B(112)) xor (A(75) and B(111)) xor (A(76) and B(110)) xor (A(77) and B(109)) xor (A(78) and B(108)) xor (A(79) and B(107)) xor (A(80) and B(106)) xor (A(81) and B(105)) xor (A(82) and B(104)) xor (A(83) and B(103)) xor (A(84) and B(102)) xor (A(85) and B(101)) xor (A(86) and B(100)) xor (A(87) and B(99)) xor (A(88) and B(98)) xor (A(89) and B(97)) xor (A(90) and B(96)) xor (A(91) and B(95)) xor (A(92) and B(94)) xor (A(93) and B(93)) xor (A(94) and B(92)) xor (A(95) and B(91)) xor (A(96) and B(90)) xor (A(97) and B(89)) xor (A(98) and B(88)) xor (A(99) and B(87)) xor (A(100) and B(86)) xor (A(101) and B(85)) xor (A(102) and B(84)) xor (A(103) and B(83)) xor (A(104) and B(82)) xor (A(105) and B(81)) xor (A(106) and B(80)) xor (A(107) and B(79)) xor (A(108) and B(78)) xor (A(109) and B(77)) xor (A(110) and B(76)) xor (A(111) and B(75)) xor (A(112) and B(74)) xor (A(113) and B(73)) xor (A(114) and B(72)) xor (A(115) and B(71)) xor (A(116) and B(70)) xor (A(117) and B(69)) xor (A(118) and B(68)) xor (A(119) and B(67)) xor (A(120) and B(66)) xor (A(121) and B(65)) xor (A(122) and B(64)) xor (A(123) and B(63)) xor (A(124) and B(62)) xor (A(125) and B(61)) xor (A(126) and B(61));
    C(60)  <= (A(0) and B(60)) xor (A(1) and B(59)) xor (A(2) and B(58)) xor (A(3) and B(57)) xor (A(4) and B(56)) xor (A(5) and B(55)) xor (A(6) and B(54)) xor (A(7) and B(53)) xor (A(8) and B(52)) xor (A(9) and B(51)) xor (A(10) and B(50)) xor (A(11) and B(49)) xor (A(12) and B(48)) xor (A(13) and B(47)) xor (A(14) and B(46)) xor (A(15) and B(45)) xor (A(16) and B(44)) xor (A(17) and B(43)) xor (A(18) and B(42)) xor (A(19) and B(41)) xor (A(20) and B(40)) xor (A(21) and B(39)) xor (A(23) and B(38)) xor (A(23) and B(37)) xor (A(24) and B(36)) xor (A(25) and B(35)) xor (A(26) and B(34)) xor (A(27) and B(33)) xor (A(28) and B(32)) xor (A(29) and B(31)) xor (A(30) and B(30)) xor (A(31) and B(29)) xor (A(32) and B(28)) xor (A(33) and B(27)) xor (A(34) and B(26)) xor (A(35) and B(25)) xor (A(36) and B(24)) xor (A(37) and B(23)) xor (A(38) and B(23)) xor (A(39) and B(21)) xor (A(40) and B(20)) xor (A(41) and B(19)) xor (A(42) and B(18)) xor (A(43) and B(17)) xor (A(44) and B(16)) xor (A(45) and B(15)) xor (A(46) and B(14)) xor (A(47) and B(13)) xor (A(48) and B(12)) xor (A(49) and B(11)) xor (A(50) and B(10)) xor (A(51) and B(9)) xor (A(52) and B(8)) xor (A(53) and B(7)) xor (A(54) and B(6)) xor (A(55) and B(5)) xor (A(56) and B(4)) xor (A(57) and B(3)) xor (A(58) and B(2)) xor (A(59) and B(1)) xor (A(60) and B(0)) xor (A(53) and B(127)) xor (A(54) and B(126)) xor (A(55) and B(125)) xor (A(56) and B(124)) xor (A(57) and B(123)) xor (A(58) and B(122)) xor (A(59) and B(121)) xor (A(60) and B(120)) xor (A(61) and B(119)) xor (A(62) and B(118)) xor (A(63) and B(117)) xor (A(64) and B(116)) xor (A(65) and B(115)) xor (A(66) and B(114)) xor (A(67) and B(113)) xor (A(68) and B(112)) xor (A(69) and B(111)) xor (A(70) and B(110)) xor (A(71) and B(109)) xor (A(72) and B(108)) xor (A(73) and B(107)) xor (A(74) and B(106)) xor (A(75) and B(105)) xor (A(76) and B(104)) xor (A(77) and B(103)) xor (A(78) and B(102)) xor (A(79) and B(101)) xor (A(80) and B(100)) xor (A(81) and B(99)) xor (A(82) and B(98)) xor (A(83) and B(97)) xor (A(84) and B(96)) xor (A(85) and B(95)) xor (A(86) and B(94)) xor (A(87) and B(93)) xor (A(88) and B(92)) xor (A(89) and B(91)) xor (A(90) and B(90)) xor (A(91) and B(89)) xor (A(92) and B(88)) xor (A(93) and B(87)) xor (A(94) and B(86)) xor (A(95) and B(85)) xor (A(96) and B(84)) xor (A(97) and B(83)) xor (A(98) and B(82)) xor (A(99) and B(81)) xor (A(100) and B(80)) xor (A(101) and B(79)) xor (A(102) and B(78)) xor (A(103) and B(77)) xor (A(104) and B(76)) xor (A(105) and B(75)) xor (A(106) and B(74)) xor (A(107) and B(73)) xor (A(108) and B(72)) xor (A(109) and B(71)) xor (A(110) and B(70)) xor (A(111) and B(69)) xor (A(112) and B(68)) xor (A(113) and B(67)) xor (A(114) and B(66)) xor (A(115) and B(65)) xor (A(116) and B(64)) xor (A(117) and B(63)) xor (A(118) and B(62)) xor (A(119) and B(61)) xor (A(120) and B(60)) xor (A(121) and B(59)) xor (A(122) and B(58)) xor (A(123) and B(57)) xor (A(124) and B(56)) xor (A(125) and B(55)) xor (A(126) and B(54)) xor (A(58) and B(127)) xor (A(59) and B(126)) xor (A(60) and B(125)) xor (A(61) and B(124)) xor (A(62) and B(123)) xor (A(63) and B(122)) xor (A(64) and B(121)) xor (A(65) and B(120)) xor (A(66) and B(119)) xor (A(67) and B(118)) xor (A(68) and B(117)) xor (A(69) and B(116)) xor (A(70) and B(115)) xor (A(71) and B(114)) xor (A(72) and B(113)) xor (A(73) and B(112)) xor (A(74) and B(111)) xor (A(75) and B(110)) xor (A(76) and B(109)) xor (A(77) and B(108)) xor (A(78) and B(107)) xor (A(79) and B(106)) xor (A(80) and B(105)) xor (A(81) and B(104)) xor (A(82) and B(103)) xor (A(83) and B(102)) xor (A(84) and B(101)) xor (A(85) and B(100)) xor (A(86) and B(99)) xor (A(87) and B(98)) xor (A(88) and B(97)) xor (A(89) and B(96)) xor (A(90) and B(95)) xor (A(91) and B(94)) xor (A(92) and B(93)) xor (A(93) and B(92)) xor (A(94) and B(91)) xor (A(95) and B(90)) xor (A(96) and B(89)) xor (A(97) and B(88)) xor (A(98) and B(87)) xor (A(99) and B(86)) xor (A(100) and B(85)) xor (A(101) and B(84)) xor (A(102) and B(83)) xor (A(103) and B(82)) xor (A(104) and B(81)) xor (A(105) and B(80)) xor (A(106) and B(79)) xor (A(107) and B(78)) xor (A(108) and B(77)) xor (A(109) and B(76)) xor (A(110) and B(75)) xor (A(111) and B(74)) xor (A(112) and B(73)) xor (A(113) and B(72)) xor (A(114) and B(71)) xor (A(115) and B(70)) xor (A(116) and B(69)) xor (A(117) and B(68)) xor (A(118) and B(67)) xor (A(119) and B(66)) xor (A(120) and B(65)) xor (A(121) and B(64)) xor (A(122) and B(63)) xor (A(123) and B(62)) xor (A(124) and B(61)) xor (A(125) and B(60)) xor (A(126) and B(59)) xor (A(59) and B(127)) xor (A(60) and B(126)) xor (A(61) and B(125)) xor (A(62) and B(124)) xor (A(63) and B(123)) xor (A(64) and B(122)) xor (A(65) and B(121)) xor (A(66) and B(120)) xor (A(67) and B(119)) xor (A(68) and B(118)) xor (A(69) and B(117)) xor (A(70) and B(116)) xor (A(71) and B(115)) xor (A(72) and B(114)) xor (A(73) and B(113)) xor (A(74) and B(112)) xor (A(75) and B(111)) xor (A(76) and B(110)) xor (A(77) and B(109)) xor (A(78) and B(108)) xor (A(79) and B(107)) xor (A(80) and B(106)) xor (A(81) and B(105)) xor (A(82) and B(104)) xor (A(83) and B(103)) xor (A(84) and B(102)) xor (A(85) and B(101)) xor (A(86) and B(100)) xor (A(87) and B(99)) xor (A(88) and B(98)) xor (A(89) and B(97)) xor (A(90) and B(96)) xor (A(91) and B(95)) xor (A(92) and B(94)) xor (A(93) and B(93)) xor (A(94) and B(92)) xor (A(95) and B(91)) xor (A(96) and B(90)) xor (A(97) and B(89)) xor (A(98) and B(88)) xor (A(99) and B(87)) xor (A(100) and B(86)) xor (A(101) and B(85)) xor (A(102) and B(84)) xor (A(103) and B(83)) xor (A(104) and B(82)) xor (A(105) and B(81)) xor (A(106) and B(80)) xor (A(107) and B(79)) xor (A(108) and B(78)) xor (A(109) and B(77)) xor (A(110) and B(76)) xor (A(111) and B(75)) xor (A(112) and B(74)) xor (A(113) and B(73)) xor (A(114) and B(72)) xor (A(115) and B(71)) xor (A(116) and B(70)) xor (A(117) and B(69)) xor (A(118) and B(68)) xor (A(119) and B(67)) xor (A(120) and B(66)) xor (A(121) and B(65)) xor (A(122) and B(64)) xor (A(123) and B(63)) xor (A(124) and B(62)) xor (A(125) and B(61)) xor (A(126) and B(60)) xor (A(60) and B(127)) xor (A(61) and B(126)) xor (A(62) and B(125)) xor (A(63) and B(124)) xor (A(64) and B(123)) xor (A(65) and B(122)) xor (A(66) and B(121)) xor (A(67) and B(120)) xor (A(68) and B(119)) xor (A(69) and B(118)) xor (A(70) and B(117)) xor (A(71) and B(116)) xor (A(72) and B(115)) xor (A(73) and B(114)) xor (A(74) and B(113)) xor (A(75) and B(112)) xor (A(76) and B(111)) xor (A(77) and B(110)) xor (A(78) and B(109)) xor (A(79) and B(108)) xor (A(80) and B(107)) xor (A(81) and B(106)) xor (A(82) and B(105)) xor (A(83) and B(104)) xor (A(84) and B(103)) xor (A(85) and B(102)) xor (A(86) and B(101)) xor (A(87) and B(100)) xor (A(88) and B(99)) xor (A(89) and B(98)) xor (A(90) and B(97)) xor (A(91) and B(96)) xor (A(92) and B(95)) xor (A(93) and B(94)) xor (A(94) and B(93)) xor (A(95) and B(92)) xor (A(96) and B(91)) xor (A(97) and B(90)) xor (A(98) and B(89)) xor (A(99) and B(88)) xor (A(100) and B(87)) xor (A(101) and B(86)) xor (A(102) and B(85)) xor (A(103) and B(84)) xor (A(104) and B(83)) xor (A(105) and B(82)) xor (A(106) and B(81)) xor (A(107) and B(80)) xor (A(108) and B(79)) xor (A(109) and B(78)) xor (A(110) and B(77)) xor (A(111) and B(76)) xor (A(112) and B(75)) xor (A(113) and B(74)) xor (A(114) and B(73)) xor (A(115) and B(72)) xor (A(116) and B(71)) xor (A(117) and B(70)) xor (A(118) and B(69)) xor (A(119) and B(68)) xor (A(120) and B(67)) xor (A(121) and B(66)) xor (A(122) and B(65)) xor (A(123) and B(64)) xor (A(124) and B(63)) xor (A(125) and B(62)) xor (A(126) and B(62));
    C(61)  <= (A(0) and B(61)) xor (A(1) and B(60)) xor (A(2) and B(59)) xor (A(3) and B(58)) xor (A(4) and B(57)) xor (A(5) and B(56)) xor (A(6) and B(55)) xor (A(7) and B(54)) xor (A(8) and B(53)) xor (A(9) and B(52)) xor (A(10) and B(51)) xor (A(11) and B(50)) xor (A(12) and B(49)) xor (A(13) and B(48)) xor (A(14) and B(47)) xor (A(15) and B(46)) xor (A(16) and B(45)) xor (A(17) and B(44)) xor (A(18) and B(43)) xor (A(19) and B(42)) xor (A(20) and B(41)) xor (A(21) and B(40)) xor (A(23) and B(39)) xor (A(23) and B(38)) xor (A(24) and B(37)) xor (A(25) and B(36)) xor (A(26) and B(35)) xor (A(27) and B(34)) xor (A(28) and B(33)) xor (A(29) and B(32)) xor (A(30) and B(31)) xor (A(31) and B(30)) xor (A(32) and B(29)) xor (A(33) and B(28)) xor (A(34) and B(27)) xor (A(35) and B(26)) xor (A(36) and B(25)) xor (A(37) and B(24)) xor (A(38) and B(23)) xor (A(39) and B(23)) xor (A(40) and B(21)) xor (A(41) and B(20)) xor (A(42) and B(19)) xor (A(43) and B(18)) xor (A(44) and B(17)) xor (A(45) and B(16)) xor (A(46) and B(15)) xor (A(47) and B(14)) xor (A(48) and B(13)) xor (A(49) and B(12)) xor (A(50) and B(11)) xor (A(51) and B(10)) xor (A(52) and B(9)) xor (A(53) and B(8)) xor (A(54) and B(7)) xor (A(55) and B(6)) xor (A(56) and B(5)) xor (A(57) and B(4)) xor (A(58) and B(3)) xor (A(59) and B(2)) xor (A(60) and B(1)) xor (A(61) and B(0)) xor (A(54) and B(127)) xor (A(55) and B(126)) xor (A(56) and B(125)) xor (A(57) and B(124)) xor (A(58) and B(123)) xor (A(59) and B(122)) xor (A(60) and B(121)) xor (A(61) and B(120)) xor (A(62) and B(119)) xor (A(63) and B(118)) xor (A(64) and B(117)) xor (A(65) and B(116)) xor (A(66) and B(115)) xor (A(67) and B(114)) xor (A(68) and B(113)) xor (A(69) and B(112)) xor (A(70) and B(111)) xor (A(71) and B(110)) xor (A(72) and B(109)) xor (A(73) and B(108)) xor (A(74) and B(107)) xor (A(75) and B(106)) xor (A(76) and B(105)) xor (A(77) and B(104)) xor (A(78) and B(103)) xor (A(79) and B(102)) xor (A(80) and B(101)) xor (A(81) and B(100)) xor (A(82) and B(99)) xor (A(83) and B(98)) xor (A(84) and B(97)) xor (A(85) and B(96)) xor (A(86) and B(95)) xor (A(87) and B(94)) xor (A(88) and B(93)) xor (A(89) and B(92)) xor (A(90) and B(91)) xor (A(91) and B(90)) xor (A(92) and B(89)) xor (A(93) and B(88)) xor (A(94) and B(87)) xor (A(95) and B(86)) xor (A(96) and B(85)) xor (A(97) and B(84)) xor (A(98) and B(83)) xor (A(99) and B(82)) xor (A(100) and B(81)) xor (A(101) and B(80)) xor (A(102) and B(79)) xor (A(103) and B(78)) xor (A(104) and B(77)) xor (A(105) and B(76)) xor (A(106) and B(75)) xor (A(107) and B(74)) xor (A(108) and B(73)) xor (A(109) and B(72)) xor (A(110) and B(71)) xor (A(111) and B(70)) xor (A(112) and B(69)) xor (A(113) and B(68)) xor (A(114) and B(67)) xor (A(115) and B(66)) xor (A(116) and B(65)) xor (A(117) and B(64)) xor (A(118) and B(63)) xor (A(119) and B(62)) xor (A(120) and B(61)) xor (A(121) and B(60)) xor (A(122) and B(59)) xor (A(123) and B(58)) xor (A(124) and B(57)) xor (A(125) and B(56)) xor (A(126) and B(55)) xor (A(59) and B(127)) xor (A(60) and B(126)) xor (A(61) and B(125)) xor (A(62) and B(124)) xor (A(63) and B(123)) xor (A(64) and B(122)) xor (A(65) and B(121)) xor (A(66) and B(120)) xor (A(67) and B(119)) xor (A(68) and B(118)) xor (A(69) and B(117)) xor (A(70) and B(116)) xor (A(71) and B(115)) xor (A(72) and B(114)) xor (A(73) and B(113)) xor (A(74) and B(112)) xor (A(75) and B(111)) xor (A(76) and B(110)) xor (A(77) and B(109)) xor (A(78) and B(108)) xor (A(79) and B(107)) xor (A(80) and B(106)) xor (A(81) and B(105)) xor (A(82) and B(104)) xor (A(83) and B(103)) xor (A(84) and B(102)) xor (A(85) and B(101)) xor (A(86) and B(100)) xor (A(87) and B(99)) xor (A(88) and B(98)) xor (A(89) and B(97)) xor (A(90) and B(96)) xor (A(91) and B(95)) xor (A(92) and B(94)) xor (A(93) and B(93)) xor (A(94) and B(92)) xor (A(95) and B(91)) xor (A(96) and B(90)) xor (A(97) and B(89)) xor (A(98) and B(88)) xor (A(99) and B(87)) xor (A(100) and B(86)) xor (A(101) and B(85)) xor (A(102) and B(84)) xor (A(103) and B(83)) xor (A(104) and B(82)) xor (A(105) and B(81)) xor (A(106) and B(80)) xor (A(107) and B(79)) xor (A(108) and B(78)) xor (A(109) and B(77)) xor (A(110) and B(76)) xor (A(111) and B(75)) xor (A(112) and B(74)) xor (A(113) and B(73)) xor (A(114) and B(72)) xor (A(115) and B(71)) xor (A(116) and B(70)) xor (A(117) and B(69)) xor (A(118) and B(68)) xor (A(119) and B(67)) xor (A(120) and B(66)) xor (A(121) and B(65)) xor (A(122) and B(64)) xor (A(123) and B(63)) xor (A(124) and B(62)) xor (A(125) and B(61)) xor (A(126) and B(60)) xor (A(60) and B(127)) xor (A(61) and B(126)) xor (A(62) and B(125)) xor (A(63) and B(124)) xor (A(64) and B(123)) xor (A(65) and B(122)) xor (A(66) and B(121)) xor (A(67) and B(120)) xor (A(68) and B(119)) xor (A(69) and B(118)) xor (A(70) and B(117)) xor (A(71) and B(116)) xor (A(72) and B(115)) xor (A(73) and B(114)) xor (A(74) and B(113)) xor (A(75) and B(112)) xor (A(76) and B(111)) xor (A(77) and B(110)) xor (A(78) and B(109)) xor (A(79) and B(108)) xor (A(80) and B(107)) xor (A(81) and B(106)) xor (A(82) and B(105)) xor (A(83) and B(104)) xor (A(84) and B(103)) xor (A(85) and B(102)) xor (A(86) and B(101)) xor (A(87) and B(100)) xor (A(88) and B(99)) xor (A(89) and B(98)) xor (A(90) and B(97)) xor (A(91) and B(96)) xor (A(92) and B(95)) xor (A(93) and B(94)) xor (A(94) and B(93)) xor (A(95) and B(92)) xor (A(96) and B(91)) xor (A(97) and B(90)) xor (A(98) and B(89)) xor (A(99) and B(88)) xor (A(100) and B(87)) xor (A(101) and B(86)) xor (A(102) and B(85)) xor (A(103) and B(84)) xor (A(104) and B(83)) xor (A(105) and B(82)) xor (A(106) and B(81)) xor (A(107) and B(80)) xor (A(108) and B(79)) xor (A(109) and B(78)) xor (A(110) and B(77)) xor (A(111) and B(76)) xor (A(112) and B(75)) xor (A(113) and B(74)) xor (A(114) and B(73)) xor (A(115) and B(72)) xor (A(116) and B(71)) xor (A(117) and B(70)) xor (A(118) and B(69)) xor (A(119) and B(68)) xor (A(120) and B(67)) xor (A(121) and B(66)) xor (A(122) and B(65)) xor (A(123) and B(64)) xor (A(124) and B(63)) xor (A(125) and B(62)) xor (A(126) and B(61)) xor (A(61) and B(127)) xor (A(62) and B(126)) xor (A(63) and B(125)) xor (A(64) and B(124)) xor (A(65) and B(123)) xor (A(66) and B(122)) xor (A(67) and B(121)) xor (A(68) and B(120)) xor (A(69) and B(119)) xor (A(70) and B(118)) xor (A(71) and B(117)) xor (A(72) and B(116)) xor (A(73) and B(115)) xor (A(74) and B(114)) xor (A(75) and B(113)) xor (A(76) and B(112)) xor (A(77) and B(111)) xor (A(78) and B(110)) xor (A(79) and B(109)) xor (A(80) and B(108)) xor (A(81) and B(107)) xor (A(82) and B(106)) xor (A(83) and B(105)) xor (A(84) and B(104)) xor (A(85) and B(103)) xor (A(86) and B(102)) xor (A(87) and B(101)) xor (A(88) and B(100)) xor (A(89) and B(99)) xor (A(90) and B(98)) xor (A(91) and B(97)) xor (A(92) and B(96)) xor (A(93) and B(95)) xor (A(94) and B(94)) xor (A(95) and B(93)) xor (A(96) and B(92)) xor (A(97) and B(91)) xor (A(98) and B(90)) xor (A(99) and B(89)) xor (A(100) and B(88)) xor (A(101) and B(87)) xor (A(102) and B(86)) xor (A(103) and B(85)) xor (A(104) and B(84)) xor (A(105) and B(83)) xor (A(106) and B(82)) xor (A(107) and B(81)) xor (A(108) and B(80)) xor (A(109) and B(79)) xor (A(110) and B(78)) xor (A(111) and B(77)) xor (A(112) and B(76)) xor (A(113) and B(75)) xor (A(114) and B(74)) xor (A(115) and B(73)) xor (A(116) and B(72)) xor (A(117) and B(71)) xor (A(118) and B(70)) xor (A(119) and B(69)) xor (A(120) and B(68)) xor (A(121) and B(67)) xor (A(122) and B(66)) xor (A(123) and B(65)) xor (A(124) and B(64)) xor (A(125) and B(63)) xor (A(126) and B(63));
    C(62)  <= (A(0) and B(62)) xor (A(1) and B(61)) xor (A(2) and B(60)) xor (A(3) and B(59)) xor (A(4) and B(58)) xor (A(5) and B(57)) xor (A(6) and B(56)) xor (A(7) and B(55)) xor (A(8) and B(54)) xor (A(9) and B(53)) xor (A(10) and B(52)) xor (A(11) and B(51)) xor (A(12) and B(50)) xor (A(13) and B(49)) xor (A(14) and B(48)) xor (A(15) and B(47)) xor (A(16) and B(46)) xor (A(17) and B(45)) xor (A(18) and B(44)) xor (A(19) and B(43)) xor (A(20) and B(42)) xor (A(21) and B(41)) xor (A(23) and B(40)) xor (A(23) and B(39)) xor (A(24) and B(38)) xor (A(25) and B(37)) xor (A(26) and B(36)) xor (A(27) and B(35)) xor (A(28) and B(34)) xor (A(29) and B(33)) xor (A(30) and B(32)) xor (A(31) and B(31)) xor (A(32) and B(30)) xor (A(33) and B(29)) xor (A(34) and B(28)) xor (A(35) and B(27)) xor (A(36) and B(26)) xor (A(37) and B(25)) xor (A(38) and B(24)) xor (A(39) and B(23)) xor (A(40) and B(23)) xor (A(41) and B(21)) xor (A(42) and B(20)) xor (A(43) and B(19)) xor (A(44) and B(18)) xor (A(45) and B(17)) xor (A(46) and B(16)) xor (A(47) and B(15)) xor (A(48) and B(14)) xor (A(49) and B(13)) xor (A(50) and B(12)) xor (A(51) and B(11)) xor (A(52) and B(10)) xor (A(53) and B(9)) xor (A(54) and B(8)) xor (A(55) and B(7)) xor (A(56) and B(6)) xor (A(57) and B(5)) xor (A(58) and B(4)) xor (A(59) and B(3)) xor (A(60) and B(2)) xor (A(61) and B(1)) xor (A(62) and B(0)) xor (A(55) and B(127)) xor (A(56) and B(126)) xor (A(57) and B(125)) xor (A(58) and B(124)) xor (A(59) and B(123)) xor (A(60) and B(122)) xor (A(61) and B(121)) xor (A(62) and B(120)) xor (A(63) and B(119)) xor (A(64) and B(118)) xor (A(65) and B(117)) xor (A(66) and B(116)) xor (A(67) and B(115)) xor (A(68) and B(114)) xor (A(69) and B(113)) xor (A(70) and B(112)) xor (A(71) and B(111)) xor (A(72) and B(110)) xor (A(73) and B(109)) xor (A(74) and B(108)) xor (A(75) and B(107)) xor (A(76) and B(106)) xor (A(77) and B(105)) xor (A(78) and B(104)) xor (A(79) and B(103)) xor (A(80) and B(102)) xor (A(81) and B(101)) xor (A(82) and B(100)) xor (A(83) and B(99)) xor (A(84) and B(98)) xor (A(85) and B(97)) xor (A(86) and B(96)) xor (A(87) and B(95)) xor (A(88) and B(94)) xor (A(89) and B(93)) xor (A(90) and B(92)) xor (A(91) and B(91)) xor (A(92) and B(90)) xor (A(93) and B(89)) xor (A(94) and B(88)) xor (A(95) and B(87)) xor (A(96) and B(86)) xor (A(97) and B(85)) xor (A(98) and B(84)) xor (A(99) and B(83)) xor (A(100) and B(82)) xor (A(101) and B(81)) xor (A(102) and B(80)) xor (A(103) and B(79)) xor (A(104) and B(78)) xor (A(105) and B(77)) xor (A(106) and B(76)) xor (A(107) and B(75)) xor (A(108) and B(74)) xor (A(109) and B(73)) xor (A(110) and B(72)) xor (A(111) and B(71)) xor (A(112) and B(70)) xor (A(113) and B(69)) xor (A(114) and B(68)) xor (A(115) and B(67)) xor (A(116) and B(66)) xor (A(117) and B(65)) xor (A(118) and B(64)) xor (A(119) and B(63)) xor (A(120) and B(62)) xor (A(121) and B(61)) xor (A(122) and B(60)) xor (A(123) and B(59)) xor (A(124) and B(58)) xor (A(125) and B(57)) xor (A(126) and B(56)) xor (A(60) and B(127)) xor (A(61) and B(126)) xor (A(62) and B(125)) xor (A(63) and B(124)) xor (A(64) and B(123)) xor (A(65) and B(122)) xor (A(66) and B(121)) xor (A(67) and B(120)) xor (A(68) and B(119)) xor (A(69) and B(118)) xor (A(70) and B(117)) xor (A(71) and B(116)) xor (A(72) and B(115)) xor (A(73) and B(114)) xor (A(74) and B(113)) xor (A(75) and B(112)) xor (A(76) and B(111)) xor (A(77) and B(110)) xor (A(78) and B(109)) xor (A(79) and B(108)) xor (A(80) and B(107)) xor (A(81) and B(106)) xor (A(82) and B(105)) xor (A(83) and B(104)) xor (A(84) and B(103)) xor (A(85) and B(102)) xor (A(86) and B(101)) xor (A(87) and B(100)) xor (A(88) and B(99)) xor (A(89) and B(98)) xor (A(90) and B(97)) xor (A(91) and B(96)) xor (A(92) and B(95)) xor (A(93) and B(94)) xor (A(94) and B(93)) xor (A(95) and B(92)) xor (A(96) and B(91)) xor (A(97) and B(90)) xor (A(98) and B(89)) xor (A(99) and B(88)) xor (A(100) and B(87)) xor (A(101) and B(86)) xor (A(102) and B(85)) xor (A(103) and B(84)) xor (A(104) and B(83)) xor (A(105) and B(82)) xor (A(106) and B(81)) xor (A(107) and B(80)) xor (A(108) and B(79)) xor (A(109) and B(78)) xor (A(110) and B(77)) xor (A(111) and B(76)) xor (A(112) and B(75)) xor (A(113) and B(74)) xor (A(114) and B(73)) xor (A(115) and B(72)) xor (A(116) and B(71)) xor (A(117) and B(70)) xor (A(118) and B(69)) xor (A(119) and B(68)) xor (A(120) and B(67)) xor (A(121) and B(66)) xor (A(122) and B(65)) xor (A(123) and B(64)) xor (A(124) and B(63)) xor (A(125) and B(62)) xor (A(126) and B(61)) xor (A(61) and B(127)) xor (A(62) and B(126)) xor (A(63) and B(125)) xor (A(64) and B(124)) xor (A(65) and B(123)) xor (A(66) and B(122)) xor (A(67) and B(121)) xor (A(68) and B(120)) xor (A(69) and B(119)) xor (A(70) and B(118)) xor (A(71) and B(117)) xor (A(72) and B(116)) xor (A(73) and B(115)) xor (A(74) and B(114)) xor (A(75) and B(113)) xor (A(76) and B(112)) xor (A(77) and B(111)) xor (A(78) and B(110)) xor (A(79) and B(109)) xor (A(80) and B(108)) xor (A(81) and B(107)) xor (A(82) and B(106)) xor (A(83) and B(105)) xor (A(84) and B(104)) xor (A(85) and B(103)) xor (A(86) and B(102)) xor (A(87) and B(101)) xor (A(88) and B(100)) xor (A(89) and B(99)) xor (A(90) and B(98)) xor (A(91) and B(97)) xor (A(92) and B(96)) xor (A(93) and B(95)) xor (A(94) and B(94)) xor (A(95) and B(93)) xor (A(96) and B(92)) xor (A(97) and B(91)) xor (A(98) and B(90)) xor (A(99) and B(89)) xor (A(100) and B(88)) xor (A(101) and B(87)) xor (A(102) and B(86)) xor (A(103) and B(85)) xor (A(104) and B(84)) xor (A(105) and B(83)) xor (A(106) and B(82)) xor (A(107) and B(81)) xor (A(108) and B(80)) xor (A(109) and B(79)) xor (A(110) and B(78)) xor (A(111) and B(77)) xor (A(112) and B(76)) xor (A(113) and B(75)) xor (A(114) and B(74)) xor (A(115) and B(73)) xor (A(116) and B(72)) xor (A(117) and B(71)) xor (A(118) and B(70)) xor (A(119) and B(69)) xor (A(120) and B(68)) xor (A(121) and B(67)) xor (A(122) and B(66)) xor (A(123) and B(65)) xor (A(124) and B(64)) xor (A(125) and B(63)) xor (A(126) and B(62)) xor (A(62) and B(127)) xor (A(63) and B(126)) xor (A(64) and B(125)) xor (A(65) and B(124)) xor (A(66) and B(123)) xor (A(67) and B(122)) xor (A(68) and B(121)) xor (A(69) and B(120)) xor (A(70) and B(119)) xor (A(71) and B(118)) xor (A(72) and B(117)) xor (A(73) and B(116)) xor (A(74) and B(115)) xor (A(75) and B(114)) xor (A(76) and B(113)) xor (A(77) and B(112)) xor (A(78) and B(111)) xor (A(79) and B(110)) xor (A(80) and B(109)) xor (A(81) and B(108)) xor (A(82) and B(107)) xor (A(83) and B(106)) xor (A(84) and B(105)) xor (A(85) and B(104)) xor (A(86) and B(103)) xor (A(87) and B(102)) xor (A(88) and B(101)) xor (A(89) and B(100)) xor (A(90) and B(99)) xor (A(91) and B(98)) xor (A(92) and B(97)) xor (A(93) and B(96)) xor (A(94) and B(95)) xor (A(95) and B(94)) xor (A(96) and B(93)) xor (A(97) and B(92)) xor (A(98) and B(91)) xor (A(99) and B(90)) xor (A(100) and B(89)) xor (A(101) and B(88)) xor (A(102) and B(87)) xor (A(103) and B(86)) xor (A(104) and B(85)) xor (A(105) and B(84)) xor (A(106) and B(83)) xor (A(107) and B(82)) xor (A(108) and B(81)) xor (A(109) and B(80)) xor (A(110) and B(79)) xor (A(111) and B(78)) xor (A(112) and B(77)) xor (A(113) and B(76)) xor (A(114) and B(75)) xor (A(115) and B(74)) xor (A(116) and B(73)) xor (A(117) and B(72)) xor (A(118) and B(71)) xor (A(119) and B(70)) xor (A(120) and B(69)) xor (A(121) and B(68)) xor (A(122) and B(67)) xor (A(123) and B(66)) xor (A(124) and B(65)) xor (A(125) and B(64)) xor (A(126) and B(64));
    C(63)  <= (A(0) and B(63)) xor (A(1) and B(62)) xor (A(2) and B(61)) xor (A(3) and B(60)) xor (A(4) and B(59)) xor (A(5) and B(58)) xor (A(6) and B(57)) xor (A(7) and B(56)) xor (A(8) and B(55)) xor (A(9) and B(54)) xor (A(10) and B(53)) xor (A(11) and B(52)) xor (A(12) and B(51)) xor (A(13) and B(50)) xor (A(14) and B(49)) xor (A(15) and B(48)) xor (A(16) and B(47)) xor (A(17) and B(46)) xor (A(18) and B(45)) xor (A(19) and B(44)) xor (A(20) and B(43)) xor (A(21) and B(42)) xor (A(23) and B(41)) xor (A(23) and B(40)) xor (A(24) and B(39)) xor (A(25) and B(38)) xor (A(26) and B(37)) xor (A(27) and B(36)) xor (A(28) and B(35)) xor (A(29) and B(34)) xor (A(30) and B(33)) xor (A(31) and B(32)) xor (A(32) and B(31)) xor (A(33) and B(30)) xor (A(34) and B(29)) xor (A(35) and B(28)) xor (A(36) and B(27)) xor (A(37) and B(26)) xor (A(38) and B(25)) xor (A(39) and B(24)) xor (A(40) and B(23)) xor (A(41) and B(23)) xor (A(42) and B(21)) xor (A(43) and B(20)) xor (A(44) and B(19)) xor (A(45) and B(18)) xor (A(46) and B(17)) xor (A(47) and B(16)) xor (A(48) and B(15)) xor (A(49) and B(14)) xor (A(50) and B(13)) xor (A(51) and B(12)) xor (A(52) and B(11)) xor (A(53) and B(10)) xor (A(54) and B(9)) xor (A(55) and B(8)) xor (A(56) and B(7)) xor (A(57) and B(6)) xor (A(58) and B(5)) xor (A(59) and B(4)) xor (A(60) and B(3)) xor (A(61) and B(2)) xor (A(62) and B(1)) xor (A(63) and B(0)) xor (A(56) and B(127)) xor (A(57) and B(126)) xor (A(58) and B(125)) xor (A(59) and B(124)) xor (A(60) and B(123)) xor (A(61) and B(122)) xor (A(62) and B(121)) xor (A(63) and B(120)) xor (A(64) and B(119)) xor (A(65) and B(118)) xor (A(66) and B(117)) xor (A(67) and B(116)) xor (A(68) and B(115)) xor (A(69) and B(114)) xor (A(70) and B(113)) xor (A(71) and B(112)) xor (A(72) and B(111)) xor (A(73) and B(110)) xor (A(74) and B(109)) xor (A(75) and B(108)) xor (A(76) and B(107)) xor (A(77) and B(106)) xor (A(78) and B(105)) xor (A(79) and B(104)) xor (A(80) and B(103)) xor (A(81) and B(102)) xor (A(82) and B(101)) xor (A(83) and B(100)) xor (A(84) and B(99)) xor (A(85) and B(98)) xor (A(86) and B(97)) xor (A(87) and B(96)) xor (A(88) and B(95)) xor (A(89) and B(94)) xor (A(90) and B(93)) xor (A(91) and B(92)) xor (A(92) and B(91)) xor (A(93) and B(90)) xor (A(94) and B(89)) xor (A(95) and B(88)) xor (A(96) and B(87)) xor (A(97) and B(86)) xor (A(98) and B(85)) xor (A(99) and B(84)) xor (A(100) and B(83)) xor (A(101) and B(82)) xor (A(102) and B(81)) xor (A(103) and B(80)) xor (A(104) and B(79)) xor (A(105) and B(78)) xor (A(106) and B(77)) xor (A(107) and B(76)) xor (A(108) and B(75)) xor (A(109) and B(74)) xor (A(110) and B(73)) xor (A(111) and B(72)) xor (A(112) and B(71)) xor (A(113) and B(70)) xor (A(114) and B(69)) xor (A(115) and B(68)) xor (A(116) and B(67)) xor (A(117) and B(66)) xor (A(118) and B(65)) xor (A(119) and B(64)) xor (A(120) and B(63)) xor (A(121) and B(62)) xor (A(122) and B(61)) xor (A(123) and B(60)) xor (A(124) and B(59)) xor (A(125) and B(58)) xor (A(126) and B(57)) xor (A(61) and B(127)) xor (A(62) and B(126)) xor (A(63) and B(125)) xor (A(64) and B(124)) xor (A(65) and B(123)) xor (A(66) and B(122)) xor (A(67) and B(121)) xor (A(68) and B(120)) xor (A(69) and B(119)) xor (A(70) and B(118)) xor (A(71) and B(117)) xor (A(72) and B(116)) xor (A(73) and B(115)) xor (A(74) and B(114)) xor (A(75) and B(113)) xor (A(76) and B(112)) xor (A(77) and B(111)) xor (A(78) and B(110)) xor (A(79) and B(109)) xor (A(80) and B(108)) xor (A(81) and B(107)) xor (A(82) and B(106)) xor (A(83) and B(105)) xor (A(84) and B(104)) xor (A(85) and B(103)) xor (A(86) and B(102)) xor (A(87) and B(101)) xor (A(88) and B(100)) xor (A(89) and B(99)) xor (A(90) and B(98)) xor (A(91) and B(97)) xor (A(92) and B(96)) xor (A(93) and B(95)) xor (A(94) and B(94)) xor (A(95) and B(93)) xor (A(96) and B(92)) xor (A(97) and B(91)) xor (A(98) and B(90)) xor (A(99) and B(89)) xor (A(100) and B(88)) xor (A(101) and B(87)) xor (A(102) and B(86)) xor (A(103) and B(85)) xor (A(104) and B(84)) xor (A(105) and B(83)) xor (A(106) and B(82)) xor (A(107) and B(81)) xor (A(108) and B(80)) xor (A(109) and B(79)) xor (A(110) and B(78)) xor (A(111) and B(77)) xor (A(112) and B(76)) xor (A(113) and B(75)) xor (A(114) and B(74)) xor (A(115) and B(73)) xor (A(116) and B(72)) xor (A(117) and B(71)) xor (A(118) and B(70)) xor (A(119) and B(69)) xor (A(120) and B(68)) xor (A(121) and B(67)) xor (A(122) and B(66)) xor (A(123) and B(65)) xor (A(124) and B(64)) xor (A(125) and B(63)) xor (A(126) and B(62)) xor (A(62) and B(127)) xor (A(63) and B(126)) xor (A(64) and B(125)) xor (A(65) and B(124)) xor (A(66) and B(123)) xor (A(67) and B(122)) xor (A(68) and B(121)) xor (A(69) and B(120)) xor (A(70) and B(119)) xor (A(71) and B(118)) xor (A(72) and B(117)) xor (A(73) and B(116)) xor (A(74) and B(115)) xor (A(75) and B(114)) xor (A(76) and B(113)) xor (A(77) and B(112)) xor (A(78) and B(111)) xor (A(79) and B(110)) xor (A(80) and B(109)) xor (A(81) and B(108)) xor (A(82) and B(107)) xor (A(83) and B(106)) xor (A(84) and B(105)) xor (A(85) and B(104)) xor (A(86) and B(103)) xor (A(87) and B(102)) xor (A(88) and B(101)) xor (A(89) and B(100)) xor (A(90) and B(99)) xor (A(91) and B(98)) xor (A(92) and B(97)) xor (A(93) and B(96)) xor (A(94) and B(95)) xor (A(95) and B(94)) xor (A(96) and B(93)) xor (A(97) and B(92)) xor (A(98) and B(91)) xor (A(99) and B(90)) xor (A(100) and B(89)) xor (A(101) and B(88)) xor (A(102) and B(87)) xor (A(103) and B(86)) xor (A(104) and B(85)) xor (A(105) and B(84)) xor (A(106) and B(83)) xor (A(107) and B(82)) xor (A(108) and B(81)) xor (A(109) and B(80)) xor (A(110) and B(79)) xor (A(111) and B(78)) xor (A(112) and B(77)) xor (A(113) and B(76)) xor (A(114) and B(75)) xor (A(115) and B(74)) xor (A(116) and B(73)) xor (A(117) and B(72)) xor (A(118) and B(71)) xor (A(119) and B(70)) xor (A(120) and B(69)) xor (A(121) and B(68)) xor (A(122) and B(67)) xor (A(123) and B(66)) xor (A(124) and B(65)) xor (A(125) and B(64)) xor (A(126) and B(63)) xor (A(63) and B(127)) xor (A(64) and B(126)) xor (A(65) and B(125)) xor (A(66) and B(124)) xor (A(67) and B(123)) xor (A(68) and B(122)) xor (A(69) and B(121)) xor (A(70) and B(120)) xor (A(71) and B(119)) xor (A(72) and B(118)) xor (A(73) and B(117)) xor (A(74) and B(116)) xor (A(75) and B(115)) xor (A(76) and B(114)) xor (A(77) and B(113)) xor (A(78) and B(112)) xor (A(79) and B(111)) xor (A(80) and B(110)) xor (A(81) and B(109)) xor (A(82) and B(108)) xor (A(83) and B(107)) xor (A(84) and B(106)) xor (A(85) and B(105)) xor (A(86) and B(104)) xor (A(87) and B(103)) xor (A(88) and B(102)) xor (A(89) and B(101)) xor (A(90) and B(100)) xor (A(91) and B(99)) xor (A(92) and B(98)) xor (A(93) and B(97)) xor (A(94) and B(96)) xor (A(95) and B(95)) xor (A(96) and B(94)) xor (A(97) and B(93)) xor (A(98) and B(92)) xor (A(99) and B(91)) xor (A(100) and B(90)) xor (A(101) and B(89)) xor (A(102) and B(88)) xor (A(103) and B(87)) xor (A(104) and B(86)) xor (A(105) and B(85)) xor (A(106) and B(84)) xor (A(107) and B(83)) xor (A(108) and B(82)) xor (A(109) and B(81)) xor (A(110) and B(80)) xor (A(111) and B(79)) xor (A(112) and B(78)) xor (A(113) and B(77)) xor (A(114) and B(76)) xor (A(115) and B(75)) xor (A(116) and B(74)) xor (A(117) and B(73)) xor (A(118) and B(72)) xor (A(119) and B(71)) xor (A(120) and B(70)) xor (A(121) and B(69)) xor (A(122) and B(68)) xor (A(123) and B(67)) xor (A(124) and B(66)) xor (A(125) and B(65)) xor (A(126) and B(65));
    C(64)  <= (A(0) and B(64)) xor (A(1) and B(63)) xor (A(2) and B(62)) xor (A(3) and B(61)) xor (A(4) and B(60)) xor (A(5) and B(59)) xor (A(6) and B(58)) xor (A(7) and B(57)) xor (A(8) and B(56)) xor (A(9) and B(55)) xor (A(10) and B(54)) xor (A(11) and B(53)) xor (A(12) and B(52)) xor (A(13) and B(51)) xor (A(14) and B(50)) xor (A(15) and B(49)) xor (A(16) and B(48)) xor (A(17) and B(47)) xor (A(18) and B(46)) xor (A(19) and B(45)) xor (A(20) and B(44)) xor (A(21) and B(43)) xor (A(23) and B(42)) xor (A(23) and B(41)) xor (A(24) and B(40)) xor (A(25) and B(39)) xor (A(26) and B(38)) xor (A(27) and B(37)) xor (A(28) and B(36)) xor (A(29) and B(35)) xor (A(30) and B(34)) xor (A(31) and B(33)) xor (A(32) and B(32)) xor (A(33) and B(31)) xor (A(34) and B(30)) xor (A(35) and B(29)) xor (A(36) and B(28)) xor (A(37) and B(27)) xor (A(38) and B(26)) xor (A(39) and B(25)) xor (A(40) and B(24)) xor (A(41) and B(23)) xor (A(42) and B(23)) xor (A(43) and B(21)) xor (A(44) and B(20)) xor (A(45) and B(19)) xor (A(46) and B(18)) xor (A(47) and B(17)) xor (A(48) and B(16)) xor (A(49) and B(15)) xor (A(50) and B(14)) xor (A(51) and B(13)) xor (A(52) and B(12)) xor (A(53) and B(11)) xor (A(54) and B(10)) xor (A(55) and B(9)) xor (A(56) and B(8)) xor (A(57) and B(7)) xor (A(58) and B(6)) xor (A(59) and B(5)) xor (A(60) and B(4)) xor (A(61) and B(3)) xor (A(62) and B(2)) xor (A(63) and B(1)) xor (A(64) and B(0)) xor (A(57) and B(127)) xor (A(58) and B(126)) xor (A(59) and B(125)) xor (A(60) and B(124)) xor (A(61) and B(123)) xor (A(62) and B(122)) xor (A(63) and B(121)) xor (A(64) and B(120)) xor (A(65) and B(119)) xor (A(66) and B(118)) xor (A(67) and B(117)) xor (A(68) and B(116)) xor (A(69) and B(115)) xor (A(70) and B(114)) xor (A(71) and B(113)) xor (A(72) and B(112)) xor (A(73) and B(111)) xor (A(74) and B(110)) xor (A(75) and B(109)) xor (A(76) and B(108)) xor (A(77) and B(107)) xor (A(78) and B(106)) xor (A(79) and B(105)) xor (A(80) and B(104)) xor (A(81) and B(103)) xor (A(82) and B(102)) xor (A(83) and B(101)) xor (A(84) and B(100)) xor (A(85) and B(99)) xor (A(86) and B(98)) xor (A(87) and B(97)) xor (A(88) and B(96)) xor (A(89) and B(95)) xor (A(90) and B(94)) xor (A(91) and B(93)) xor (A(92) and B(92)) xor (A(93) and B(91)) xor (A(94) and B(90)) xor (A(95) and B(89)) xor (A(96) and B(88)) xor (A(97) and B(87)) xor (A(98) and B(86)) xor (A(99) and B(85)) xor (A(100) and B(84)) xor (A(101) and B(83)) xor (A(102) and B(82)) xor (A(103) and B(81)) xor (A(104) and B(80)) xor (A(105) and B(79)) xor (A(106) and B(78)) xor (A(107) and B(77)) xor (A(108) and B(76)) xor (A(109) and B(75)) xor (A(110) and B(74)) xor (A(111) and B(73)) xor (A(112) and B(72)) xor (A(113) and B(71)) xor (A(114) and B(70)) xor (A(115) and B(69)) xor (A(116) and B(68)) xor (A(117) and B(67)) xor (A(118) and B(66)) xor (A(119) and B(65)) xor (A(120) and B(64)) xor (A(121) and B(63)) xor (A(122) and B(62)) xor (A(123) and B(61)) xor (A(124) and B(60)) xor (A(125) and B(59)) xor (A(126) and B(58)) xor (A(62) and B(127)) xor (A(63) and B(126)) xor (A(64) and B(125)) xor (A(65) and B(124)) xor (A(66) and B(123)) xor (A(67) and B(122)) xor (A(68) and B(121)) xor (A(69) and B(120)) xor (A(70) and B(119)) xor (A(71) and B(118)) xor (A(72) and B(117)) xor (A(73) and B(116)) xor (A(74) and B(115)) xor (A(75) and B(114)) xor (A(76) and B(113)) xor (A(77) and B(112)) xor (A(78) and B(111)) xor (A(79) and B(110)) xor (A(80) and B(109)) xor (A(81) and B(108)) xor (A(82) and B(107)) xor (A(83) and B(106)) xor (A(84) and B(105)) xor (A(85) and B(104)) xor (A(86) and B(103)) xor (A(87) and B(102)) xor (A(88) and B(101)) xor (A(89) and B(100)) xor (A(90) and B(99)) xor (A(91) and B(98)) xor (A(92) and B(97)) xor (A(93) and B(96)) xor (A(94) and B(95)) xor (A(95) and B(94)) xor (A(96) and B(93)) xor (A(97) and B(92)) xor (A(98) and B(91)) xor (A(99) and B(90)) xor (A(100) and B(89)) xor (A(101) and B(88)) xor (A(102) and B(87)) xor (A(103) and B(86)) xor (A(104) and B(85)) xor (A(105) and B(84)) xor (A(106) and B(83)) xor (A(107) and B(82)) xor (A(108) and B(81)) xor (A(109) and B(80)) xor (A(110) and B(79)) xor (A(111) and B(78)) xor (A(112) and B(77)) xor (A(113) and B(76)) xor (A(114) and B(75)) xor (A(115) and B(74)) xor (A(116) and B(73)) xor (A(117) and B(72)) xor (A(118) and B(71)) xor (A(119) and B(70)) xor (A(120) and B(69)) xor (A(121) and B(68)) xor (A(122) and B(67)) xor (A(123) and B(66)) xor (A(124) and B(65)) xor (A(125) and B(64)) xor (A(126) and B(63)) xor (A(63) and B(127)) xor (A(64) and B(126)) xor (A(65) and B(125)) xor (A(66) and B(124)) xor (A(67) and B(123)) xor (A(68) and B(122)) xor (A(69) and B(121)) xor (A(70) and B(120)) xor (A(71) and B(119)) xor (A(72) and B(118)) xor (A(73) and B(117)) xor (A(74) and B(116)) xor (A(75) and B(115)) xor (A(76) and B(114)) xor (A(77) and B(113)) xor (A(78) and B(112)) xor (A(79) and B(111)) xor (A(80) and B(110)) xor (A(81) and B(109)) xor (A(82) and B(108)) xor (A(83) and B(107)) xor (A(84) and B(106)) xor (A(85) and B(105)) xor (A(86) and B(104)) xor (A(87) and B(103)) xor (A(88) and B(102)) xor (A(89) and B(101)) xor (A(90) and B(100)) xor (A(91) and B(99)) xor (A(92) and B(98)) xor (A(93) and B(97)) xor (A(94) and B(96)) xor (A(95) and B(95)) xor (A(96) and B(94)) xor (A(97) and B(93)) xor (A(98) and B(92)) xor (A(99) and B(91)) xor (A(100) and B(90)) xor (A(101) and B(89)) xor (A(102) and B(88)) xor (A(103) and B(87)) xor (A(104) and B(86)) xor (A(105) and B(85)) xor (A(106) and B(84)) xor (A(107) and B(83)) xor (A(108) and B(82)) xor (A(109) and B(81)) xor (A(110) and B(80)) xor (A(111) and B(79)) xor (A(112) and B(78)) xor (A(113) and B(77)) xor (A(114) and B(76)) xor (A(115) and B(75)) xor (A(116) and B(74)) xor (A(117) and B(73)) xor (A(118) and B(72)) xor (A(119) and B(71)) xor (A(120) and B(70)) xor (A(121) and B(69)) xor (A(122) and B(68)) xor (A(123) and B(67)) xor (A(124) and B(66)) xor (A(125) and B(65)) xor (A(126) and B(64)) xor (A(64) and B(127)) xor (A(65) and B(126)) xor (A(66) and B(125)) xor (A(67) and B(124)) xor (A(68) and B(123)) xor (A(69) and B(122)) xor (A(70) and B(121)) xor (A(71) and B(120)) xor (A(72) and B(119)) xor (A(73) and B(118)) xor (A(74) and B(117)) xor (A(75) and B(116)) xor (A(76) and B(115)) xor (A(77) and B(114)) xor (A(78) and B(113)) xor (A(79) and B(112)) xor (A(80) and B(111)) xor (A(81) and B(110)) xor (A(82) and B(109)) xor (A(83) and B(108)) xor (A(84) and B(107)) xor (A(85) and B(106)) xor (A(86) and B(105)) xor (A(87) and B(104)) xor (A(88) and B(103)) xor (A(89) and B(102)) xor (A(90) and B(101)) xor (A(91) and B(100)) xor (A(92) and B(99)) xor (A(93) and B(98)) xor (A(94) and B(97)) xor (A(95) and B(96)) xor (A(96) and B(95)) xor (A(97) and B(94)) xor (A(98) and B(93)) xor (A(99) and B(92)) xor (A(100) and B(91)) xor (A(101) and B(90)) xor (A(102) and B(89)) xor (A(103) and B(88)) xor (A(104) and B(87)) xor (A(105) and B(86)) xor (A(106) and B(85)) xor (A(107) and B(84)) xor (A(108) and B(83)) xor (A(109) and B(82)) xor (A(110) and B(81)) xor (A(111) and B(80)) xor (A(112) and B(79)) xor (A(113) and B(78)) xor (A(114) and B(77)) xor (A(115) and B(76)) xor (A(116) and B(75)) xor (A(117) and B(74)) xor (A(118) and B(73)) xor (A(119) and B(72)) xor (A(120) and B(71)) xor (A(121) and B(70)) xor (A(122) and B(69)) xor (A(123) and B(68)) xor (A(124) and B(67)) xor (A(125) and B(66)) xor (A(126) and B(66));
    C(65)  <= (A(0) and B(65)) xor (A(1) and B(64)) xor (A(2) and B(63)) xor (A(3) and B(62)) xor (A(4) and B(61)) xor (A(5) and B(60)) xor (A(6) and B(59)) xor (A(7) and B(58)) xor (A(8) and B(57)) xor (A(9) and B(56)) xor (A(10) and B(55)) xor (A(11) and B(54)) xor (A(12) and B(53)) xor (A(13) and B(52)) xor (A(14) and B(51)) xor (A(15) and B(50)) xor (A(16) and B(49)) xor (A(17) and B(48)) xor (A(18) and B(47)) xor (A(19) and B(46)) xor (A(20) and B(45)) xor (A(21) and B(44)) xor (A(23) and B(43)) xor (A(23) and B(42)) xor (A(24) and B(41)) xor (A(25) and B(40)) xor (A(26) and B(39)) xor (A(27) and B(38)) xor (A(28) and B(37)) xor (A(29) and B(36)) xor (A(30) and B(35)) xor (A(31) and B(34)) xor (A(32) and B(33)) xor (A(33) and B(32)) xor (A(34) and B(31)) xor (A(35) and B(30)) xor (A(36) and B(29)) xor (A(37) and B(28)) xor (A(38) and B(27)) xor (A(39) and B(26)) xor (A(40) and B(25)) xor (A(41) and B(24)) xor (A(42) and B(23)) xor (A(43) and B(23)) xor (A(44) and B(21)) xor (A(45) and B(20)) xor (A(46) and B(19)) xor (A(47) and B(18)) xor (A(48) and B(17)) xor (A(49) and B(16)) xor (A(50) and B(15)) xor (A(51) and B(14)) xor (A(52) and B(13)) xor (A(53) and B(12)) xor (A(54) and B(11)) xor (A(55) and B(10)) xor (A(56) and B(9)) xor (A(57) and B(8)) xor (A(58) and B(7)) xor (A(59) and B(6)) xor (A(60) and B(5)) xor (A(61) and B(4)) xor (A(62) and B(3)) xor (A(63) and B(2)) xor (A(64) and B(1)) xor (A(65) and B(0)) xor (A(58) and B(127)) xor (A(59) and B(126)) xor (A(60) and B(125)) xor (A(61) and B(124)) xor (A(62) and B(123)) xor (A(63) and B(122)) xor (A(64) and B(121)) xor (A(65) and B(120)) xor (A(66) and B(119)) xor (A(67) and B(118)) xor (A(68) and B(117)) xor (A(69) and B(116)) xor (A(70) and B(115)) xor (A(71) and B(114)) xor (A(72) and B(113)) xor (A(73) and B(112)) xor (A(74) and B(111)) xor (A(75) and B(110)) xor (A(76) and B(109)) xor (A(77) and B(108)) xor (A(78) and B(107)) xor (A(79) and B(106)) xor (A(80) and B(105)) xor (A(81) and B(104)) xor (A(82) and B(103)) xor (A(83) and B(102)) xor (A(84) and B(101)) xor (A(85) and B(100)) xor (A(86) and B(99)) xor (A(87) and B(98)) xor (A(88) and B(97)) xor (A(89) and B(96)) xor (A(90) and B(95)) xor (A(91) and B(94)) xor (A(92) and B(93)) xor (A(93) and B(92)) xor (A(94) and B(91)) xor (A(95) and B(90)) xor (A(96) and B(89)) xor (A(97) and B(88)) xor (A(98) and B(87)) xor (A(99) and B(86)) xor (A(100) and B(85)) xor (A(101) and B(84)) xor (A(102) and B(83)) xor (A(103) and B(82)) xor (A(104) and B(81)) xor (A(105) and B(80)) xor (A(106) and B(79)) xor (A(107) and B(78)) xor (A(108) and B(77)) xor (A(109) and B(76)) xor (A(110) and B(75)) xor (A(111) and B(74)) xor (A(112) and B(73)) xor (A(113) and B(72)) xor (A(114) and B(71)) xor (A(115) and B(70)) xor (A(116) and B(69)) xor (A(117) and B(68)) xor (A(118) and B(67)) xor (A(119) and B(66)) xor (A(120) and B(65)) xor (A(121) and B(64)) xor (A(122) and B(63)) xor (A(123) and B(62)) xor (A(124) and B(61)) xor (A(125) and B(60)) xor (A(126) and B(59)) xor (A(63) and B(127)) xor (A(64) and B(126)) xor (A(65) and B(125)) xor (A(66) and B(124)) xor (A(67) and B(123)) xor (A(68) and B(122)) xor (A(69) and B(121)) xor (A(70) and B(120)) xor (A(71) and B(119)) xor (A(72) and B(118)) xor (A(73) and B(117)) xor (A(74) and B(116)) xor (A(75) and B(115)) xor (A(76) and B(114)) xor (A(77) and B(113)) xor (A(78) and B(112)) xor (A(79) and B(111)) xor (A(80) and B(110)) xor (A(81) and B(109)) xor (A(82) and B(108)) xor (A(83) and B(107)) xor (A(84) and B(106)) xor (A(85) and B(105)) xor (A(86) and B(104)) xor (A(87) and B(103)) xor (A(88) and B(102)) xor (A(89) and B(101)) xor (A(90) and B(100)) xor (A(91) and B(99)) xor (A(92) and B(98)) xor (A(93) and B(97)) xor (A(94) and B(96)) xor (A(95) and B(95)) xor (A(96) and B(94)) xor (A(97) and B(93)) xor (A(98) and B(92)) xor (A(99) and B(91)) xor (A(100) and B(90)) xor (A(101) and B(89)) xor (A(102) and B(88)) xor (A(103) and B(87)) xor (A(104) and B(86)) xor (A(105) and B(85)) xor (A(106) and B(84)) xor (A(107) and B(83)) xor (A(108) and B(82)) xor (A(109) and B(81)) xor (A(110) and B(80)) xor (A(111) and B(79)) xor (A(112) and B(78)) xor (A(113) and B(77)) xor (A(114) and B(76)) xor (A(115) and B(75)) xor (A(116) and B(74)) xor (A(117) and B(73)) xor (A(118) and B(72)) xor (A(119) and B(71)) xor (A(120) and B(70)) xor (A(121) and B(69)) xor (A(122) and B(68)) xor (A(123) and B(67)) xor (A(124) and B(66)) xor (A(125) and B(65)) xor (A(126) and B(64)) xor (A(64) and B(127)) xor (A(65) and B(126)) xor (A(66) and B(125)) xor (A(67) and B(124)) xor (A(68) and B(123)) xor (A(69) and B(122)) xor (A(70) and B(121)) xor (A(71) and B(120)) xor (A(72) and B(119)) xor (A(73) and B(118)) xor (A(74) and B(117)) xor (A(75) and B(116)) xor (A(76) and B(115)) xor (A(77) and B(114)) xor (A(78) and B(113)) xor (A(79) and B(112)) xor (A(80) and B(111)) xor (A(81) and B(110)) xor (A(82) and B(109)) xor (A(83) and B(108)) xor (A(84) and B(107)) xor (A(85) and B(106)) xor (A(86) and B(105)) xor (A(87) and B(104)) xor (A(88) and B(103)) xor (A(89) and B(102)) xor (A(90) and B(101)) xor (A(91) and B(100)) xor (A(92) and B(99)) xor (A(93) and B(98)) xor (A(94) and B(97)) xor (A(95) and B(96)) xor (A(96) and B(95)) xor (A(97) and B(94)) xor (A(98) and B(93)) xor (A(99) and B(92)) xor (A(100) and B(91)) xor (A(101) and B(90)) xor (A(102) and B(89)) xor (A(103) and B(88)) xor (A(104) and B(87)) xor (A(105) and B(86)) xor (A(106) and B(85)) xor (A(107) and B(84)) xor (A(108) and B(83)) xor (A(109) and B(82)) xor (A(110) and B(81)) xor (A(111) and B(80)) xor (A(112) and B(79)) xor (A(113) and B(78)) xor (A(114) and B(77)) xor (A(115) and B(76)) xor (A(116) and B(75)) xor (A(117) and B(74)) xor (A(118) and B(73)) xor (A(119) and B(72)) xor (A(120) and B(71)) xor (A(121) and B(70)) xor (A(122) and B(69)) xor (A(123) and B(68)) xor (A(124) and B(67)) xor (A(125) and B(66)) xor (A(126) and B(65)) xor (A(65) and B(127)) xor (A(66) and B(126)) xor (A(67) and B(125)) xor (A(68) and B(124)) xor (A(69) and B(123)) xor (A(70) and B(122)) xor (A(71) and B(121)) xor (A(72) and B(120)) xor (A(73) and B(119)) xor (A(74) and B(118)) xor (A(75) and B(117)) xor (A(76) and B(116)) xor (A(77) and B(115)) xor (A(78) and B(114)) xor (A(79) and B(113)) xor (A(80) and B(112)) xor (A(81) and B(111)) xor (A(82) and B(110)) xor (A(83) and B(109)) xor (A(84) and B(108)) xor (A(85) and B(107)) xor (A(86) and B(106)) xor (A(87) and B(105)) xor (A(88) and B(104)) xor (A(89) and B(103)) xor (A(90) and B(102)) xor (A(91) and B(101)) xor (A(92) and B(100)) xor (A(93) and B(99)) xor (A(94) and B(98)) xor (A(95) and B(97)) xor (A(96) and B(96)) xor (A(97) and B(95)) xor (A(98) and B(94)) xor (A(99) and B(93)) xor (A(100) and B(92)) xor (A(101) and B(91)) xor (A(102) and B(90)) xor (A(103) and B(89)) xor (A(104) and B(88)) xor (A(105) and B(87)) xor (A(106) and B(86)) xor (A(107) and B(85)) xor (A(108) and B(84)) xor (A(109) and B(83)) xor (A(110) and B(82)) xor (A(111) and B(81)) xor (A(112) and B(80)) xor (A(113) and B(79)) xor (A(114) and B(78)) xor (A(115) and B(77)) xor (A(116) and B(76)) xor (A(117) and B(75)) xor (A(118) and B(74)) xor (A(119) and B(73)) xor (A(120) and B(72)) xor (A(121) and B(71)) xor (A(122) and B(70)) xor (A(123) and B(69)) xor (A(124) and B(68)) xor (A(125) and B(67)) xor (A(126) and B(67));
    C(66)  <= (A(0) and B(66)) xor (A(1) and B(65)) xor (A(2) and B(64)) xor (A(3) and B(63)) xor (A(4) and B(62)) xor (A(5) and B(61)) xor (A(6) and B(60)) xor (A(7) and B(59)) xor (A(8) and B(58)) xor (A(9) and B(57)) xor (A(10) and B(56)) xor (A(11) and B(55)) xor (A(12) and B(54)) xor (A(13) and B(53)) xor (A(14) and B(52)) xor (A(15) and B(51)) xor (A(16) and B(50)) xor (A(17) and B(49)) xor (A(18) and B(48)) xor (A(19) and B(47)) xor (A(20) and B(46)) xor (A(21) and B(45)) xor (A(23) and B(44)) xor (A(23) and B(43)) xor (A(24) and B(42)) xor (A(25) and B(41)) xor (A(26) and B(40)) xor (A(27) and B(39)) xor (A(28) and B(38)) xor (A(29) and B(37)) xor (A(30) and B(36)) xor (A(31) and B(35)) xor (A(32) and B(34)) xor (A(33) and B(33)) xor (A(34) and B(32)) xor (A(35) and B(31)) xor (A(36) and B(30)) xor (A(37) and B(29)) xor (A(38) and B(28)) xor (A(39) and B(27)) xor (A(40) and B(26)) xor (A(41) and B(25)) xor (A(42) and B(24)) xor (A(43) and B(23)) xor (A(44) and B(23)) xor (A(45) and B(21)) xor (A(46) and B(20)) xor (A(47) and B(19)) xor (A(48) and B(18)) xor (A(49) and B(17)) xor (A(50) and B(16)) xor (A(51) and B(15)) xor (A(52) and B(14)) xor (A(53) and B(13)) xor (A(54) and B(12)) xor (A(55) and B(11)) xor (A(56) and B(10)) xor (A(57) and B(9)) xor (A(58) and B(8)) xor (A(59) and B(7)) xor (A(60) and B(6)) xor (A(61) and B(5)) xor (A(62) and B(4)) xor (A(63) and B(3)) xor (A(64) and B(2)) xor (A(65) and B(1)) xor (A(66) and B(0)) xor (A(59) and B(127)) xor (A(60) and B(126)) xor (A(61) and B(125)) xor (A(62) and B(124)) xor (A(63) and B(123)) xor (A(64) and B(122)) xor (A(65) and B(121)) xor (A(66) and B(120)) xor (A(67) and B(119)) xor (A(68) and B(118)) xor (A(69) and B(117)) xor (A(70) and B(116)) xor (A(71) and B(115)) xor (A(72) and B(114)) xor (A(73) and B(113)) xor (A(74) and B(112)) xor (A(75) and B(111)) xor (A(76) and B(110)) xor (A(77) and B(109)) xor (A(78) and B(108)) xor (A(79) and B(107)) xor (A(80) and B(106)) xor (A(81) and B(105)) xor (A(82) and B(104)) xor (A(83) and B(103)) xor (A(84) and B(102)) xor (A(85) and B(101)) xor (A(86) and B(100)) xor (A(87) and B(99)) xor (A(88) and B(98)) xor (A(89) and B(97)) xor (A(90) and B(96)) xor (A(91) and B(95)) xor (A(92) and B(94)) xor (A(93) and B(93)) xor (A(94) and B(92)) xor (A(95) and B(91)) xor (A(96) and B(90)) xor (A(97) and B(89)) xor (A(98) and B(88)) xor (A(99) and B(87)) xor (A(100) and B(86)) xor (A(101) and B(85)) xor (A(102) and B(84)) xor (A(103) and B(83)) xor (A(104) and B(82)) xor (A(105) and B(81)) xor (A(106) and B(80)) xor (A(107) and B(79)) xor (A(108) and B(78)) xor (A(109) and B(77)) xor (A(110) and B(76)) xor (A(111) and B(75)) xor (A(112) and B(74)) xor (A(113) and B(73)) xor (A(114) and B(72)) xor (A(115) and B(71)) xor (A(116) and B(70)) xor (A(117) and B(69)) xor (A(118) and B(68)) xor (A(119) and B(67)) xor (A(120) and B(66)) xor (A(121) and B(65)) xor (A(122) and B(64)) xor (A(123) and B(63)) xor (A(124) and B(62)) xor (A(125) and B(61)) xor (A(126) and B(60)) xor (A(64) and B(127)) xor (A(65) and B(126)) xor (A(66) and B(125)) xor (A(67) and B(124)) xor (A(68) and B(123)) xor (A(69) and B(122)) xor (A(70) and B(121)) xor (A(71) and B(120)) xor (A(72) and B(119)) xor (A(73) and B(118)) xor (A(74) and B(117)) xor (A(75) and B(116)) xor (A(76) and B(115)) xor (A(77) and B(114)) xor (A(78) and B(113)) xor (A(79) and B(112)) xor (A(80) and B(111)) xor (A(81) and B(110)) xor (A(82) and B(109)) xor (A(83) and B(108)) xor (A(84) and B(107)) xor (A(85) and B(106)) xor (A(86) and B(105)) xor (A(87) and B(104)) xor (A(88) and B(103)) xor (A(89) and B(102)) xor (A(90) and B(101)) xor (A(91) and B(100)) xor (A(92) and B(99)) xor (A(93) and B(98)) xor (A(94) and B(97)) xor (A(95) and B(96)) xor (A(96) and B(95)) xor (A(97) and B(94)) xor (A(98) and B(93)) xor (A(99) and B(92)) xor (A(100) and B(91)) xor (A(101) and B(90)) xor (A(102) and B(89)) xor (A(103) and B(88)) xor (A(104) and B(87)) xor (A(105) and B(86)) xor (A(106) and B(85)) xor (A(107) and B(84)) xor (A(108) and B(83)) xor (A(109) and B(82)) xor (A(110) and B(81)) xor (A(111) and B(80)) xor (A(112) and B(79)) xor (A(113) and B(78)) xor (A(114) and B(77)) xor (A(115) and B(76)) xor (A(116) and B(75)) xor (A(117) and B(74)) xor (A(118) and B(73)) xor (A(119) and B(72)) xor (A(120) and B(71)) xor (A(121) and B(70)) xor (A(122) and B(69)) xor (A(123) and B(68)) xor (A(124) and B(67)) xor (A(125) and B(66)) xor (A(126) and B(65)) xor (A(65) and B(127)) xor (A(66) and B(126)) xor (A(67) and B(125)) xor (A(68) and B(124)) xor (A(69) and B(123)) xor (A(70) and B(122)) xor (A(71) and B(121)) xor (A(72) and B(120)) xor (A(73) and B(119)) xor (A(74) and B(118)) xor (A(75) and B(117)) xor (A(76) and B(116)) xor (A(77) and B(115)) xor (A(78) and B(114)) xor (A(79) and B(113)) xor (A(80) and B(112)) xor (A(81) and B(111)) xor (A(82) and B(110)) xor (A(83) and B(109)) xor (A(84) and B(108)) xor (A(85) and B(107)) xor (A(86) and B(106)) xor (A(87) and B(105)) xor (A(88) and B(104)) xor (A(89) and B(103)) xor (A(90) and B(102)) xor (A(91) and B(101)) xor (A(92) and B(100)) xor (A(93) and B(99)) xor (A(94) and B(98)) xor (A(95) and B(97)) xor (A(96) and B(96)) xor (A(97) and B(95)) xor (A(98) and B(94)) xor (A(99) and B(93)) xor (A(100) and B(92)) xor (A(101) and B(91)) xor (A(102) and B(90)) xor (A(103) and B(89)) xor (A(104) and B(88)) xor (A(105) and B(87)) xor (A(106) and B(86)) xor (A(107) and B(85)) xor (A(108) and B(84)) xor (A(109) and B(83)) xor (A(110) and B(82)) xor (A(111) and B(81)) xor (A(112) and B(80)) xor (A(113) and B(79)) xor (A(114) and B(78)) xor (A(115) and B(77)) xor (A(116) and B(76)) xor (A(117) and B(75)) xor (A(118) and B(74)) xor (A(119) and B(73)) xor (A(120) and B(72)) xor (A(121) and B(71)) xor (A(122) and B(70)) xor (A(123) and B(69)) xor (A(124) and B(68)) xor (A(125) and B(67)) xor (A(126) and B(66)) xor (A(66) and B(127)) xor (A(67) and B(126)) xor (A(68) and B(125)) xor (A(69) and B(124)) xor (A(70) and B(123)) xor (A(71) and B(122)) xor (A(72) and B(121)) xor (A(73) and B(120)) xor (A(74) and B(119)) xor (A(75) and B(118)) xor (A(76) and B(117)) xor (A(77) and B(116)) xor (A(78) and B(115)) xor (A(79) and B(114)) xor (A(80) and B(113)) xor (A(81) and B(112)) xor (A(82) and B(111)) xor (A(83) and B(110)) xor (A(84) and B(109)) xor (A(85) and B(108)) xor (A(86) and B(107)) xor (A(87) and B(106)) xor (A(88) and B(105)) xor (A(89) and B(104)) xor (A(90) and B(103)) xor (A(91) and B(102)) xor (A(92) and B(101)) xor (A(93) and B(100)) xor (A(94) and B(99)) xor (A(95) and B(98)) xor (A(96) and B(97)) xor (A(97) and B(96)) xor (A(98) and B(95)) xor (A(99) and B(94)) xor (A(100) and B(93)) xor (A(101) and B(92)) xor (A(102) and B(91)) xor (A(103) and B(90)) xor (A(104) and B(89)) xor (A(105) and B(88)) xor (A(106) and B(87)) xor (A(107) and B(86)) xor (A(108) and B(85)) xor (A(109) and B(84)) xor (A(110) and B(83)) xor (A(111) and B(82)) xor (A(112) and B(81)) xor (A(113) and B(80)) xor (A(114) and B(79)) xor (A(115) and B(78)) xor (A(116) and B(77)) xor (A(117) and B(76)) xor (A(118) and B(75)) xor (A(119) and B(74)) xor (A(120) and B(73)) xor (A(121) and B(72)) xor (A(122) and B(71)) xor (A(123) and B(70)) xor (A(124) and B(69)) xor (A(125) and B(68)) xor (A(126) and B(68));
    C(67)  <= (A(0) and B(67)) xor (A(1) and B(66)) xor (A(2) and B(65)) xor (A(3) and B(64)) xor (A(4) and B(63)) xor (A(5) and B(62)) xor (A(6) and B(61)) xor (A(7) and B(60)) xor (A(8) and B(59)) xor (A(9) and B(58)) xor (A(10) and B(57)) xor (A(11) and B(56)) xor (A(12) and B(55)) xor (A(13) and B(54)) xor (A(14) and B(53)) xor (A(15) and B(52)) xor (A(16) and B(51)) xor (A(17) and B(50)) xor (A(18) and B(49)) xor (A(19) and B(48)) xor (A(20) and B(47)) xor (A(21) and B(46)) xor (A(23) and B(45)) xor (A(23) and B(44)) xor (A(24) and B(43)) xor (A(25) and B(42)) xor (A(26) and B(41)) xor (A(27) and B(40)) xor (A(28) and B(39)) xor (A(29) and B(38)) xor (A(30) and B(37)) xor (A(31) and B(36)) xor (A(32) and B(35)) xor (A(33) and B(34)) xor (A(34) and B(33)) xor (A(35) and B(32)) xor (A(36) and B(31)) xor (A(37) and B(30)) xor (A(38) and B(29)) xor (A(39) and B(28)) xor (A(40) and B(27)) xor (A(41) and B(26)) xor (A(42) and B(25)) xor (A(43) and B(24)) xor (A(44) and B(23)) xor (A(45) and B(23)) xor (A(46) and B(21)) xor (A(47) and B(20)) xor (A(48) and B(19)) xor (A(49) and B(18)) xor (A(50) and B(17)) xor (A(51) and B(16)) xor (A(52) and B(15)) xor (A(53) and B(14)) xor (A(54) and B(13)) xor (A(55) and B(12)) xor (A(56) and B(11)) xor (A(57) and B(10)) xor (A(58) and B(9)) xor (A(59) and B(8)) xor (A(60) and B(7)) xor (A(61) and B(6)) xor (A(62) and B(5)) xor (A(63) and B(4)) xor (A(64) and B(3)) xor (A(65) and B(2)) xor (A(66) and B(1)) xor (A(67) and B(0)) xor (A(60) and B(127)) xor (A(61) and B(126)) xor (A(62) and B(125)) xor (A(63) and B(124)) xor (A(64) and B(123)) xor (A(65) and B(122)) xor (A(66) and B(121)) xor (A(67) and B(120)) xor (A(68) and B(119)) xor (A(69) and B(118)) xor (A(70) and B(117)) xor (A(71) and B(116)) xor (A(72) and B(115)) xor (A(73) and B(114)) xor (A(74) and B(113)) xor (A(75) and B(112)) xor (A(76) and B(111)) xor (A(77) and B(110)) xor (A(78) and B(109)) xor (A(79) and B(108)) xor (A(80) and B(107)) xor (A(81) and B(106)) xor (A(82) and B(105)) xor (A(83) and B(104)) xor (A(84) and B(103)) xor (A(85) and B(102)) xor (A(86) and B(101)) xor (A(87) and B(100)) xor (A(88) and B(99)) xor (A(89) and B(98)) xor (A(90) and B(97)) xor (A(91) and B(96)) xor (A(92) and B(95)) xor (A(93) and B(94)) xor (A(94) and B(93)) xor (A(95) and B(92)) xor (A(96) and B(91)) xor (A(97) and B(90)) xor (A(98) and B(89)) xor (A(99) and B(88)) xor (A(100) and B(87)) xor (A(101) and B(86)) xor (A(102) and B(85)) xor (A(103) and B(84)) xor (A(104) and B(83)) xor (A(105) and B(82)) xor (A(106) and B(81)) xor (A(107) and B(80)) xor (A(108) and B(79)) xor (A(109) and B(78)) xor (A(110) and B(77)) xor (A(111) and B(76)) xor (A(112) and B(75)) xor (A(113) and B(74)) xor (A(114) and B(73)) xor (A(115) and B(72)) xor (A(116) and B(71)) xor (A(117) and B(70)) xor (A(118) and B(69)) xor (A(119) and B(68)) xor (A(120) and B(67)) xor (A(121) and B(66)) xor (A(122) and B(65)) xor (A(123) and B(64)) xor (A(124) and B(63)) xor (A(125) and B(62)) xor (A(126) and B(61)) xor (A(65) and B(127)) xor (A(66) and B(126)) xor (A(67) and B(125)) xor (A(68) and B(124)) xor (A(69) and B(123)) xor (A(70) and B(122)) xor (A(71) and B(121)) xor (A(72) and B(120)) xor (A(73) and B(119)) xor (A(74) and B(118)) xor (A(75) and B(117)) xor (A(76) and B(116)) xor (A(77) and B(115)) xor (A(78) and B(114)) xor (A(79) and B(113)) xor (A(80) and B(112)) xor (A(81) and B(111)) xor (A(82) and B(110)) xor (A(83) and B(109)) xor (A(84) and B(108)) xor (A(85) and B(107)) xor (A(86) and B(106)) xor (A(87) and B(105)) xor (A(88) and B(104)) xor (A(89) and B(103)) xor (A(90) and B(102)) xor (A(91) and B(101)) xor (A(92) and B(100)) xor (A(93) and B(99)) xor (A(94) and B(98)) xor (A(95) and B(97)) xor (A(96) and B(96)) xor (A(97) and B(95)) xor (A(98) and B(94)) xor (A(99) and B(93)) xor (A(100) and B(92)) xor (A(101) and B(91)) xor (A(102) and B(90)) xor (A(103) and B(89)) xor (A(104) and B(88)) xor (A(105) and B(87)) xor (A(106) and B(86)) xor (A(107) and B(85)) xor (A(108) and B(84)) xor (A(109) and B(83)) xor (A(110) and B(82)) xor (A(111) and B(81)) xor (A(112) and B(80)) xor (A(113) and B(79)) xor (A(114) and B(78)) xor (A(115) and B(77)) xor (A(116) and B(76)) xor (A(117) and B(75)) xor (A(118) and B(74)) xor (A(119) and B(73)) xor (A(120) and B(72)) xor (A(121) and B(71)) xor (A(122) and B(70)) xor (A(123) and B(69)) xor (A(124) and B(68)) xor (A(125) and B(67)) xor (A(126) and B(66)) xor (A(66) and B(127)) xor (A(67) and B(126)) xor (A(68) and B(125)) xor (A(69) and B(124)) xor (A(70) and B(123)) xor (A(71) and B(122)) xor (A(72) and B(121)) xor (A(73) and B(120)) xor (A(74) and B(119)) xor (A(75) and B(118)) xor (A(76) and B(117)) xor (A(77) and B(116)) xor (A(78) and B(115)) xor (A(79) and B(114)) xor (A(80) and B(113)) xor (A(81) and B(112)) xor (A(82) and B(111)) xor (A(83) and B(110)) xor (A(84) and B(109)) xor (A(85) and B(108)) xor (A(86) and B(107)) xor (A(87) and B(106)) xor (A(88) and B(105)) xor (A(89) and B(104)) xor (A(90) and B(103)) xor (A(91) and B(102)) xor (A(92) and B(101)) xor (A(93) and B(100)) xor (A(94) and B(99)) xor (A(95) and B(98)) xor (A(96) and B(97)) xor (A(97) and B(96)) xor (A(98) and B(95)) xor (A(99) and B(94)) xor (A(100) and B(93)) xor (A(101) and B(92)) xor (A(102) and B(91)) xor (A(103) and B(90)) xor (A(104) and B(89)) xor (A(105) and B(88)) xor (A(106) and B(87)) xor (A(107) and B(86)) xor (A(108) and B(85)) xor (A(109) and B(84)) xor (A(110) and B(83)) xor (A(111) and B(82)) xor (A(112) and B(81)) xor (A(113) and B(80)) xor (A(114) and B(79)) xor (A(115) and B(78)) xor (A(116) and B(77)) xor (A(117) and B(76)) xor (A(118) and B(75)) xor (A(119) and B(74)) xor (A(120) and B(73)) xor (A(121) and B(72)) xor (A(122) and B(71)) xor (A(123) and B(70)) xor (A(124) and B(69)) xor (A(125) and B(68)) xor (A(126) and B(67)) xor (A(67) and B(127)) xor (A(68) and B(126)) xor (A(69) and B(125)) xor (A(70) and B(124)) xor (A(71) and B(123)) xor (A(72) and B(122)) xor (A(73) and B(121)) xor (A(74) and B(120)) xor (A(75) and B(119)) xor (A(76) and B(118)) xor (A(77) and B(117)) xor (A(78) and B(116)) xor (A(79) and B(115)) xor (A(80) and B(114)) xor (A(81) and B(113)) xor (A(82) and B(112)) xor (A(83) and B(111)) xor (A(84) and B(110)) xor (A(85) and B(109)) xor (A(86) and B(108)) xor (A(87) and B(107)) xor (A(88) and B(106)) xor (A(89) and B(105)) xor (A(90) and B(104)) xor (A(91) and B(103)) xor (A(92) and B(102)) xor (A(93) and B(101)) xor (A(94) and B(100)) xor (A(95) and B(99)) xor (A(96) and B(98)) xor (A(97) and B(97)) xor (A(98) and B(96)) xor (A(99) and B(95)) xor (A(100) and B(94)) xor (A(101) and B(93)) xor (A(102) and B(92)) xor (A(103) and B(91)) xor (A(104) and B(90)) xor (A(105) and B(89)) xor (A(106) and B(88)) xor (A(107) and B(87)) xor (A(108) and B(86)) xor (A(109) and B(85)) xor (A(110) and B(84)) xor (A(111) and B(83)) xor (A(112) and B(82)) xor (A(113) and B(81)) xor (A(114) and B(80)) xor (A(115) and B(79)) xor (A(116) and B(78)) xor (A(117) and B(77)) xor (A(118) and B(76)) xor (A(119) and B(75)) xor (A(120) and B(74)) xor (A(121) and B(73)) xor (A(122) and B(72)) xor (A(123) and B(71)) xor (A(124) and B(70)) xor (A(125) and B(69)) xor (A(126) and B(69));
    C(68)  <= (A(0) and B(68)) xor (A(1) and B(67)) xor (A(2) and B(66)) xor (A(3) and B(65)) xor (A(4) and B(64)) xor (A(5) and B(63)) xor (A(6) and B(62)) xor (A(7) and B(61)) xor (A(8) and B(60)) xor (A(9) and B(59)) xor (A(10) and B(58)) xor (A(11) and B(57)) xor (A(12) and B(56)) xor (A(13) and B(55)) xor (A(14) and B(54)) xor (A(15) and B(53)) xor (A(16) and B(52)) xor (A(17) and B(51)) xor (A(18) and B(50)) xor (A(19) and B(49)) xor (A(20) and B(48)) xor (A(21) and B(47)) xor (A(23) and B(46)) xor (A(23) and B(45)) xor (A(24) and B(44)) xor (A(25) and B(43)) xor (A(26) and B(42)) xor (A(27) and B(41)) xor (A(28) and B(40)) xor (A(29) and B(39)) xor (A(30) and B(38)) xor (A(31) and B(37)) xor (A(32) and B(36)) xor (A(33) and B(35)) xor (A(34) and B(34)) xor (A(35) and B(33)) xor (A(36) and B(32)) xor (A(37) and B(31)) xor (A(38) and B(30)) xor (A(39) and B(29)) xor (A(40) and B(28)) xor (A(41) and B(27)) xor (A(42) and B(26)) xor (A(43) and B(25)) xor (A(44) and B(24)) xor (A(45) and B(23)) xor (A(46) and B(23)) xor (A(47) and B(21)) xor (A(48) and B(20)) xor (A(49) and B(19)) xor (A(50) and B(18)) xor (A(51) and B(17)) xor (A(52) and B(16)) xor (A(53) and B(15)) xor (A(54) and B(14)) xor (A(55) and B(13)) xor (A(56) and B(12)) xor (A(57) and B(11)) xor (A(58) and B(10)) xor (A(59) and B(9)) xor (A(60) and B(8)) xor (A(61) and B(7)) xor (A(62) and B(6)) xor (A(63) and B(5)) xor (A(64) and B(4)) xor (A(65) and B(3)) xor (A(66) and B(2)) xor (A(67) and B(1)) xor (A(68) and B(0)) xor (A(61) and B(127)) xor (A(62) and B(126)) xor (A(63) and B(125)) xor (A(64) and B(124)) xor (A(65) and B(123)) xor (A(66) and B(122)) xor (A(67) and B(121)) xor (A(68) and B(120)) xor (A(69) and B(119)) xor (A(70) and B(118)) xor (A(71) and B(117)) xor (A(72) and B(116)) xor (A(73) and B(115)) xor (A(74) and B(114)) xor (A(75) and B(113)) xor (A(76) and B(112)) xor (A(77) and B(111)) xor (A(78) and B(110)) xor (A(79) and B(109)) xor (A(80) and B(108)) xor (A(81) and B(107)) xor (A(82) and B(106)) xor (A(83) and B(105)) xor (A(84) and B(104)) xor (A(85) and B(103)) xor (A(86) and B(102)) xor (A(87) and B(101)) xor (A(88) and B(100)) xor (A(89) and B(99)) xor (A(90) and B(98)) xor (A(91) and B(97)) xor (A(92) and B(96)) xor (A(93) and B(95)) xor (A(94) and B(94)) xor (A(95) and B(93)) xor (A(96) and B(92)) xor (A(97) and B(91)) xor (A(98) and B(90)) xor (A(99) and B(89)) xor (A(100) and B(88)) xor (A(101) and B(87)) xor (A(102) and B(86)) xor (A(103) and B(85)) xor (A(104) and B(84)) xor (A(105) and B(83)) xor (A(106) and B(82)) xor (A(107) and B(81)) xor (A(108) and B(80)) xor (A(109) and B(79)) xor (A(110) and B(78)) xor (A(111) and B(77)) xor (A(112) and B(76)) xor (A(113) and B(75)) xor (A(114) and B(74)) xor (A(115) and B(73)) xor (A(116) and B(72)) xor (A(117) and B(71)) xor (A(118) and B(70)) xor (A(119) and B(69)) xor (A(120) and B(68)) xor (A(121) and B(67)) xor (A(122) and B(66)) xor (A(123) and B(65)) xor (A(124) and B(64)) xor (A(125) and B(63)) xor (A(126) and B(62)) xor (A(66) and B(127)) xor (A(67) and B(126)) xor (A(68) and B(125)) xor (A(69) and B(124)) xor (A(70) and B(123)) xor (A(71) and B(122)) xor (A(72) and B(121)) xor (A(73) and B(120)) xor (A(74) and B(119)) xor (A(75) and B(118)) xor (A(76) and B(117)) xor (A(77) and B(116)) xor (A(78) and B(115)) xor (A(79) and B(114)) xor (A(80) and B(113)) xor (A(81) and B(112)) xor (A(82) and B(111)) xor (A(83) and B(110)) xor (A(84) and B(109)) xor (A(85) and B(108)) xor (A(86) and B(107)) xor (A(87) and B(106)) xor (A(88) and B(105)) xor (A(89) and B(104)) xor (A(90) and B(103)) xor (A(91) and B(102)) xor (A(92) and B(101)) xor (A(93) and B(100)) xor (A(94) and B(99)) xor (A(95) and B(98)) xor (A(96) and B(97)) xor (A(97) and B(96)) xor (A(98) and B(95)) xor (A(99) and B(94)) xor (A(100) and B(93)) xor (A(101) and B(92)) xor (A(102) and B(91)) xor (A(103) and B(90)) xor (A(104) and B(89)) xor (A(105) and B(88)) xor (A(106) and B(87)) xor (A(107) and B(86)) xor (A(108) and B(85)) xor (A(109) and B(84)) xor (A(110) and B(83)) xor (A(111) and B(82)) xor (A(112) and B(81)) xor (A(113) and B(80)) xor (A(114) and B(79)) xor (A(115) and B(78)) xor (A(116) and B(77)) xor (A(117) and B(76)) xor (A(118) and B(75)) xor (A(119) and B(74)) xor (A(120) and B(73)) xor (A(121) and B(72)) xor (A(122) and B(71)) xor (A(123) and B(70)) xor (A(124) and B(69)) xor (A(125) and B(68)) xor (A(126) and B(67)) xor (A(67) and B(127)) xor (A(68) and B(126)) xor (A(69) and B(125)) xor (A(70) and B(124)) xor (A(71) and B(123)) xor (A(72) and B(122)) xor (A(73) and B(121)) xor (A(74) and B(120)) xor (A(75) and B(119)) xor (A(76) and B(118)) xor (A(77) and B(117)) xor (A(78) and B(116)) xor (A(79) and B(115)) xor (A(80) and B(114)) xor (A(81) and B(113)) xor (A(82) and B(112)) xor (A(83) and B(111)) xor (A(84) and B(110)) xor (A(85) and B(109)) xor (A(86) and B(108)) xor (A(87) and B(107)) xor (A(88) and B(106)) xor (A(89) and B(105)) xor (A(90) and B(104)) xor (A(91) and B(103)) xor (A(92) and B(102)) xor (A(93) and B(101)) xor (A(94) and B(100)) xor (A(95) and B(99)) xor (A(96) and B(98)) xor (A(97) and B(97)) xor (A(98) and B(96)) xor (A(99) and B(95)) xor (A(100) and B(94)) xor (A(101) and B(93)) xor (A(102) and B(92)) xor (A(103) and B(91)) xor (A(104) and B(90)) xor (A(105) and B(89)) xor (A(106) and B(88)) xor (A(107) and B(87)) xor (A(108) and B(86)) xor (A(109) and B(85)) xor (A(110) and B(84)) xor (A(111) and B(83)) xor (A(112) and B(82)) xor (A(113) and B(81)) xor (A(114) and B(80)) xor (A(115) and B(79)) xor (A(116) and B(78)) xor (A(117) and B(77)) xor (A(118) and B(76)) xor (A(119) and B(75)) xor (A(120) and B(74)) xor (A(121) and B(73)) xor (A(122) and B(72)) xor (A(123) and B(71)) xor (A(124) and B(70)) xor (A(125) and B(69)) xor (A(126) and B(68)) xor (A(68) and B(127)) xor (A(69) and B(126)) xor (A(70) and B(125)) xor (A(71) and B(124)) xor (A(72) and B(123)) xor (A(73) and B(122)) xor (A(74) and B(121)) xor (A(75) and B(120)) xor (A(76) and B(119)) xor (A(77) and B(118)) xor (A(78) and B(117)) xor (A(79) and B(116)) xor (A(80) and B(115)) xor (A(81) and B(114)) xor (A(82) and B(113)) xor (A(83) and B(112)) xor (A(84) and B(111)) xor (A(85) and B(110)) xor (A(86) and B(109)) xor (A(87) and B(108)) xor (A(88) and B(107)) xor (A(89) and B(106)) xor (A(90) and B(105)) xor (A(91) and B(104)) xor (A(92) and B(103)) xor (A(93) and B(102)) xor (A(94) and B(101)) xor (A(95) and B(100)) xor (A(96) and B(99)) xor (A(97) and B(98)) xor (A(98) and B(97)) xor (A(99) and B(96)) xor (A(100) and B(95)) xor (A(101) and B(94)) xor (A(102) and B(93)) xor (A(103) and B(92)) xor (A(104) and B(91)) xor (A(105) and B(90)) xor (A(106) and B(89)) xor (A(107) and B(88)) xor (A(108) and B(87)) xor (A(109) and B(86)) xor (A(110) and B(85)) xor (A(111) and B(84)) xor (A(112) and B(83)) xor (A(113) and B(82)) xor (A(114) and B(81)) xor (A(115) and B(80)) xor (A(116) and B(79)) xor (A(117) and B(78)) xor (A(118) and B(77)) xor (A(119) and B(76)) xor (A(120) and B(75)) xor (A(121) and B(74)) xor (A(122) and B(73)) xor (A(123) and B(72)) xor (A(124) and B(71)) xor (A(125) and B(70)) xor (A(126) and B(70));
    C(69)  <= (A(0) and B(69)) xor (A(1) and B(68)) xor (A(2) and B(67)) xor (A(3) and B(66)) xor (A(4) and B(65)) xor (A(5) and B(64)) xor (A(6) and B(63)) xor (A(7) and B(62)) xor (A(8) and B(61)) xor (A(9) and B(60)) xor (A(10) and B(59)) xor (A(11) and B(58)) xor (A(12) and B(57)) xor (A(13) and B(56)) xor (A(14) and B(55)) xor (A(15) and B(54)) xor (A(16) and B(53)) xor (A(17) and B(52)) xor (A(18) and B(51)) xor (A(19) and B(50)) xor (A(20) and B(49)) xor (A(21) and B(48)) xor (A(23) and B(47)) xor (A(23) and B(46)) xor (A(24) and B(45)) xor (A(25) and B(44)) xor (A(26) and B(43)) xor (A(27) and B(42)) xor (A(28) and B(41)) xor (A(29) and B(40)) xor (A(30) and B(39)) xor (A(31) and B(38)) xor (A(32) and B(37)) xor (A(33) and B(36)) xor (A(34) and B(35)) xor (A(35) and B(34)) xor (A(36) and B(33)) xor (A(37) and B(32)) xor (A(38) and B(31)) xor (A(39) and B(30)) xor (A(40) and B(29)) xor (A(41) and B(28)) xor (A(42) and B(27)) xor (A(43) and B(26)) xor (A(44) and B(25)) xor (A(45) and B(24)) xor (A(46) and B(23)) xor (A(47) and B(23)) xor (A(48) and B(21)) xor (A(49) and B(20)) xor (A(50) and B(19)) xor (A(51) and B(18)) xor (A(52) and B(17)) xor (A(53) and B(16)) xor (A(54) and B(15)) xor (A(55) and B(14)) xor (A(56) and B(13)) xor (A(57) and B(12)) xor (A(58) and B(11)) xor (A(59) and B(10)) xor (A(60) and B(9)) xor (A(61) and B(8)) xor (A(62) and B(7)) xor (A(63) and B(6)) xor (A(64) and B(5)) xor (A(65) and B(4)) xor (A(66) and B(3)) xor (A(67) and B(2)) xor (A(68) and B(1)) xor (A(69) and B(0)) xor (A(62) and B(127)) xor (A(63) and B(126)) xor (A(64) and B(125)) xor (A(65) and B(124)) xor (A(66) and B(123)) xor (A(67) and B(122)) xor (A(68) and B(121)) xor (A(69) and B(120)) xor (A(70) and B(119)) xor (A(71) and B(118)) xor (A(72) and B(117)) xor (A(73) and B(116)) xor (A(74) and B(115)) xor (A(75) and B(114)) xor (A(76) and B(113)) xor (A(77) and B(112)) xor (A(78) and B(111)) xor (A(79) and B(110)) xor (A(80) and B(109)) xor (A(81) and B(108)) xor (A(82) and B(107)) xor (A(83) and B(106)) xor (A(84) and B(105)) xor (A(85) and B(104)) xor (A(86) and B(103)) xor (A(87) and B(102)) xor (A(88) and B(101)) xor (A(89) and B(100)) xor (A(90) and B(99)) xor (A(91) and B(98)) xor (A(92) and B(97)) xor (A(93) and B(96)) xor (A(94) and B(95)) xor (A(95) and B(94)) xor (A(96) and B(93)) xor (A(97) and B(92)) xor (A(98) and B(91)) xor (A(99) and B(90)) xor (A(100) and B(89)) xor (A(101) and B(88)) xor (A(102) and B(87)) xor (A(103) and B(86)) xor (A(104) and B(85)) xor (A(105) and B(84)) xor (A(106) and B(83)) xor (A(107) and B(82)) xor (A(108) and B(81)) xor (A(109) and B(80)) xor (A(110) and B(79)) xor (A(111) and B(78)) xor (A(112) and B(77)) xor (A(113) and B(76)) xor (A(114) and B(75)) xor (A(115) and B(74)) xor (A(116) and B(73)) xor (A(117) and B(72)) xor (A(118) and B(71)) xor (A(119) and B(70)) xor (A(120) and B(69)) xor (A(121) and B(68)) xor (A(122) and B(67)) xor (A(123) and B(66)) xor (A(124) and B(65)) xor (A(125) and B(64)) xor (A(126) and B(63)) xor (A(67) and B(127)) xor (A(68) and B(126)) xor (A(69) and B(125)) xor (A(70) and B(124)) xor (A(71) and B(123)) xor (A(72) and B(122)) xor (A(73) and B(121)) xor (A(74) and B(120)) xor (A(75) and B(119)) xor (A(76) and B(118)) xor (A(77) and B(117)) xor (A(78) and B(116)) xor (A(79) and B(115)) xor (A(80) and B(114)) xor (A(81) and B(113)) xor (A(82) and B(112)) xor (A(83) and B(111)) xor (A(84) and B(110)) xor (A(85) and B(109)) xor (A(86) and B(108)) xor (A(87) and B(107)) xor (A(88) and B(106)) xor (A(89) and B(105)) xor (A(90) and B(104)) xor (A(91) and B(103)) xor (A(92) and B(102)) xor (A(93) and B(101)) xor (A(94) and B(100)) xor (A(95) and B(99)) xor (A(96) and B(98)) xor (A(97) and B(97)) xor (A(98) and B(96)) xor (A(99) and B(95)) xor (A(100) and B(94)) xor (A(101) and B(93)) xor (A(102) and B(92)) xor (A(103) and B(91)) xor (A(104) and B(90)) xor (A(105) and B(89)) xor (A(106) and B(88)) xor (A(107) and B(87)) xor (A(108) and B(86)) xor (A(109) and B(85)) xor (A(110) and B(84)) xor (A(111) and B(83)) xor (A(112) and B(82)) xor (A(113) and B(81)) xor (A(114) and B(80)) xor (A(115) and B(79)) xor (A(116) and B(78)) xor (A(117) and B(77)) xor (A(118) and B(76)) xor (A(119) and B(75)) xor (A(120) and B(74)) xor (A(121) and B(73)) xor (A(122) and B(72)) xor (A(123) and B(71)) xor (A(124) and B(70)) xor (A(125) and B(69)) xor (A(126) and B(68)) xor (A(68) and B(127)) xor (A(69) and B(126)) xor (A(70) and B(125)) xor (A(71) and B(124)) xor (A(72) and B(123)) xor (A(73) and B(122)) xor (A(74) and B(121)) xor (A(75) and B(120)) xor (A(76) and B(119)) xor (A(77) and B(118)) xor (A(78) and B(117)) xor (A(79) and B(116)) xor (A(80) and B(115)) xor (A(81) and B(114)) xor (A(82) and B(113)) xor (A(83) and B(112)) xor (A(84) and B(111)) xor (A(85) and B(110)) xor (A(86) and B(109)) xor (A(87) and B(108)) xor (A(88) and B(107)) xor (A(89) and B(106)) xor (A(90) and B(105)) xor (A(91) and B(104)) xor (A(92) and B(103)) xor (A(93) and B(102)) xor (A(94) and B(101)) xor (A(95) and B(100)) xor (A(96) and B(99)) xor (A(97) and B(98)) xor (A(98) and B(97)) xor (A(99) and B(96)) xor (A(100) and B(95)) xor (A(101) and B(94)) xor (A(102) and B(93)) xor (A(103) and B(92)) xor (A(104) and B(91)) xor (A(105) and B(90)) xor (A(106) and B(89)) xor (A(107) and B(88)) xor (A(108) and B(87)) xor (A(109) and B(86)) xor (A(110) and B(85)) xor (A(111) and B(84)) xor (A(112) and B(83)) xor (A(113) and B(82)) xor (A(114) and B(81)) xor (A(115) and B(80)) xor (A(116) and B(79)) xor (A(117) and B(78)) xor (A(118) and B(77)) xor (A(119) and B(76)) xor (A(120) and B(75)) xor (A(121) and B(74)) xor (A(122) and B(73)) xor (A(123) and B(72)) xor (A(124) and B(71)) xor (A(125) and B(70)) xor (A(126) and B(69)) xor (A(69) and B(127)) xor (A(70) and B(126)) xor (A(71) and B(125)) xor (A(72) and B(124)) xor (A(73) and B(123)) xor (A(74) and B(122)) xor (A(75) and B(121)) xor (A(76) and B(120)) xor (A(77) and B(119)) xor (A(78) and B(118)) xor (A(79) and B(117)) xor (A(80) and B(116)) xor (A(81) and B(115)) xor (A(82) and B(114)) xor (A(83) and B(113)) xor (A(84) and B(112)) xor (A(85) and B(111)) xor (A(86) and B(110)) xor (A(87) and B(109)) xor (A(88) and B(108)) xor (A(89) and B(107)) xor (A(90) and B(106)) xor (A(91) and B(105)) xor (A(92) and B(104)) xor (A(93) and B(103)) xor (A(94) and B(102)) xor (A(95) and B(101)) xor (A(96) and B(100)) xor (A(97) and B(99)) xor (A(98) and B(98)) xor (A(99) and B(97)) xor (A(100) and B(96)) xor (A(101) and B(95)) xor (A(102) and B(94)) xor (A(103) and B(93)) xor (A(104) and B(92)) xor (A(105) and B(91)) xor (A(106) and B(90)) xor (A(107) and B(89)) xor (A(108) and B(88)) xor (A(109) and B(87)) xor (A(110) and B(86)) xor (A(111) and B(85)) xor (A(112) and B(84)) xor (A(113) and B(83)) xor (A(114) and B(82)) xor (A(115) and B(81)) xor (A(116) and B(80)) xor (A(117) and B(79)) xor (A(118) and B(78)) xor (A(119) and B(77)) xor (A(120) and B(76)) xor (A(121) and B(75)) xor (A(122) and B(74)) xor (A(123) and B(73)) xor (A(124) and B(72)) xor (A(125) and B(71)) xor (A(126) and B(71));
    C(70)  <= (A(0) and B(70)) xor (A(1) and B(69)) xor (A(2) and B(68)) xor (A(3) and B(67)) xor (A(4) and B(66)) xor (A(5) and B(65)) xor (A(6) and B(64)) xor (A(7) and B(63)) xor (A(8) and B(62)) xor (A(9) and B(61)) xor (A(10) and B(60)) xor (A(11) and B(59)) xor (A(12) and B(58)) xor (A(13) and B(57)) xor (A(14) and B(56)) xor (A(15) and B(55)) xor (A(16) and B(54)) xor (A(17) and B(53)) xor (A(18) and B(52)) xor (A(19) and B(51)) xor (A(20) and B(50)) xor (A(21) and B(49)) xor (A(23) and B(48)) xor (A(23) and B(47)) xor (A(24) and B(46)) xor (A(25) and B(45)) xor (A(26) and B(44)) xor (A(27) and B(43)) xor (A(28) and B(42)) xor (A(29) and B(41)) xor (A(30) and B(40)) xor (A(31) and B(39)) xor (A(32) and B(38)) xor (A(33) and B(37)) xor (A(34) and B(36)) xor (A(35) and B(35)) xor (A(36) and B(34)) xor (A(37) and B(33)) xor (A(38) and B(32)) xor (A(39) and B(31)) xor (A(40) and B(30)) xor (A(41) and B(29)) xor (A(42) and B(28)) xor (A(43) and B(27)) xor (A(44) and B(26)) xor (A(45) and B(25)) xor (A(46) and B(24)) xor (A(47) and B(23)) xor (A(48) and B(23)) xor (A(49) and B(21)) xor (A(50) and B(20)) xor (A(51) and B(19)) xor (A(52) and B(18)) xor (A(53) and B(17)) xor (A(54) and B(16)) xor (A(55) and B(15)) xor (A(56) and B(14)) xor (A(57) and B(13)) xor (A(58) and B(12)) xor (A(59) and B(11)) xor (A(60) and B(10)) xor (A(61) and B(9)) xor (A(62) and B(8)) xor (A(63) and B(7)) xor (A(64) and B(6)) xor (A(65) and B(5)) xor (A(66) and B(4)) xor (A(67) and B(3)) xor (A(68) and B(2)) xor (A(69) and B(1)) xor (A(70) and B(0)) xor (A(63) and B(127)) xor (A(64) and B(126)) xor (A(65) and B(125)) xor (A(66) and B(124)) xor (A(67) and B(123)) xor (A(68) and B(122)) xor (A(69) and B(121)) xor (A(70) and B(120)) xor (A(71) and B(119)) xor (A(72) and B(118)) xor (A(73) and B(117)) xor (A(74) and B(116)) xor (A(75) and B(115)) xor (A(76) and B(114)) xor (A(77) and B(113)) xor (A(78) and B(112)) xor (A(79) and B(111)) xor (A(80) and B(110)) xor (A(81) and B(109)) xor (A(82) and B(108)) xor (A(83) and B(107)) xor (A(84) and B(106)) xor (A(85) and B(105)) xor (A(86) and B(104)) xor (A(87) and B(103)) xor (A(88) and B(102)) xor (A(89) and B(101)) xor (A(90) and B(100)) xor (A(91) and B(99)) xor (A(92) and B(98)) xor (A(93) and B(97)) xor (A(94) and B(96)) xor (A(95) and B(95)) xor (A(96) and B(94)) xor (A(97) and B(93)) xor (A(98) and B(92)) xor (A(99) and B(91)) xor (A(100) and B(90)) xor (A(101) and B(89)) xor (A(102) and B(88)) xor (A(103) and B(87)) xor (A(104) and B(86)) xor (A(105) and B(85)) xor (A(106) and B(84)) xor (A(107) and B(83)) xor (A(108) and B(82)) xor (A(109) and B(81)) xor (A(110) and B(80)) xor (A(111) and B(79)) xor (A(112) and B(78)) xor (A(113) and B(77)) xor (A(114) and B(76)) xor (A(115) and B(75)) xor (A(116) and B(74)) xor (A(117) and B(73)) xor (A(118) and B(72)) xor (A(119) and B(71)) xor (A(120) and B(70)) xor (A(121) and B(69)) xor (A(122) and B(68)) xor (A(123) and B(67)) xor (A(124) and B(66)) xor (A(125) and B(65)) xor (A(126) and B(64)) xor (A(68) and B(127)) xor (A(69) and B(126)) xor (A(70) and B(125)) xor (A(71) and B(124)) xor (A(72) and B(123)) xor (A(73) and B(122)) xor (A(74) and B(121)) xor (A(75) and B(120)) xor (A(76) and B(119)) xor (A(77) and B(118)) xor (A(78) and B(117)) xor (A(79) and B(116)) xor (A(80) and B(115)) xor (A(81) and B(114)) xor (A(82) and B(113)) xor (A(83) and B(112)) xor (A(84) and B(111)) xor (A(85) and B(110)) xor (A(86) and B(109)) xor (A(87) and B(108)) xor (A(88) and B(107)) xor (A(89) and B(106)) xor (A(90) and B(105)) xor (A(91) and B(104)) xor (A(92) and B(103)) xor (A(93) and B(102)) xor (A(94) and B(101)) xor (A(95) and B(100)) xor (A(96) and B(99)) xor (A(97) and B(98)) xor (A(98) and B(97)) xor (A(99) and B(96)) xor (A(100) and B(95)) xor (A(101) and B(94)) xor (A(102) and B(93)) xor (A(103) and B(92)) xor (A(104) and B(91)) xor (A(105) and B(90)) xor (A(106) and B(89)) xor (A(107) and B(88)) xor (A(108) and B(87)) xor (A(109) and B(86)) xor (A(110) and B(85)) xor (A(111) and B(84)) xor (A(112) and B(83)) xor (A(113) and B(82)) xor (A(114) and B(81)) xor (A(115) and B(80)) xor (A(116) and B(79)) xor (A(117) and B(78)) xor (A(118) and B(77)) xor (A(119) and B(76)) xor (A(120) and B(75)) xor (A(121) and B(74)) xor (A(122) and B(73)) xor (A(123) and B(72)) xor (A(124) and B(71)) xor (A(125) and B(70)) xor (A(126) and B(69)) xor (A(69) and B(127)) xor (A(70) and B(126)) xor (A(71) and B(125)) xor (A(72) and B(124)) xor (A(73) and B(123)) xor (A(74) and B(122)) xor (A(75) and B(121)) xor (A(76) and B(120)) xor (A(77) and B(119)) xor (A(78) and B(118)) xor (A(79) and B(117)) xor (A(80) and B(116)) xor (A(81) and B(115)) xor (A(82) and B(114)) xor (A(83) and B(113)) xor (A(84) and B(112)) xor (A(85) and B(111)) xor (A(86) and B(110)) xor (A(87) and B(109)) xor (A(88) and B(108)) xor (A(89) and B(107)) xor (A(90) and B(106)) xor (A(91) and B(105)) xor (A(92) and B(104)) xor (A(93) and B(103)) xor (A(94) and B(102)) xor (A(95) and B(101)) xor (A(96) and B(100)) xor (A(97) and B(99)) xor (A(98) and B(98)) xor (A(99) and B(97)) xor (A(100) and B(96)) xor (A(101) and B(95)) xor (A(102) and B(94)) xor (A(103) and B(93)) xor (A(104) and B(92)) xor (A(105) and B(91)) xor (A(106) and B(90)) xor (A(107) and B(89)) xor (A(108) and B(88)) xor (A(109) and B(87)) xor (A(110) and B(86)) xor (A(111) and B(85)) xor (A(112) and B(84)) xor (A(113) and B(83)) xor (A(114) and B(82)) xor (A(115) and B(81)) xor (A(116) and B(80)) xor (A(117) and B(79)) xor (A(118) and B(78)) xor (A(119) and B(77)) xor (A(120) and B(76)) xor (A(121) and B(75)) xor (A(122) and B(74)) xor (A(123) and B(73)) xor (A(124) and B(72)) xor (A(125) and B(71)) xor (A(126) and B(70)) xor (A(70) and B(127)) xor (A(71) and B(126)) xor (A(72) and B(125)) xor (A(73) and B(124)) xor (A(74) and B(123)) xor (A(75) and B(122)) xor (A(76) and B(121)) xor (A(77) and B(120)) xor (A(78) and B(119)) xor (A(79) and B(118)) xor (A(80) and B(117)) xor (A(81) and B(116)) xor (A(82) and B(115)) xor (A(83) and B(114)) xor (A(84) and B(113)) xor (A(85) and B(112)) xor (A(86) and B(111)) xor (A(87) and B(110)) xor (A(88) and B(109)) xor (A(89) and B(108)) xor (A(90) and B(107)) xor (A(91) and B(106)) xor (A(92) and B(105)) xor (A(93) and B(104)) xor (A(94) and B(103)) xor (A(95) and B(102)) xor (A(96) and B(101)) xor (A(97) and B(100)) xor (A(98) and B(99)) xor (A(99) and B(98)) xor (A(100) and B(97)) xor (A(101) and B(96)) xor (A(102) and B(95)) xor (A(103) and B(94)) xor (A(104) and B(93)) xor (A(105) and B(92)) xor (A(106) and B(91)) xor (A(107) and B(90)) xor (A(108) and B(89)) xor (A(109) and B(88)) xor (A(110) and B(87)) xor (A(111) and B(86)) xor (A(112) and B(85)) xor (A(113) and B(84)) xor (A(114) and B(83)) xor (A(115) and B(82)) xor (A(116) and B(81)) xor (A(117) and B(80)) xor (A(118) and B(79)) xor (A(119) and B(78)) xor (A(120) and B(77)) xor (A(121) and B(76)) xor (A(122) and B(75)) xor (A(123) and B(74)) xor (A(124) and B(73)) xor (A(125) and B(72)) xor (A(126) and B(72));
    C(71)  <= (A(0) and B(71)) xor (A(1) and B(70)) xor (A(2) and B(69)) xor (A(3) and B(68)) xor (A(4) and B(67)) xor (A(5) and B(66)) xor (A(6) and B(65)) xor (A(7) and B(64)) xor (A(8) and B(63)) xor (A(9) and B(62)) xor (A(10) and B(61)) xor (A(11) and B(60)) xor (A(12) and B(59)) xor (A(13) and B(58)) xor (A(14) and B(57)) xor (A(15) and B(56)) xor (A(16) and B(55)) xor (A(17) and B(54)) xor (A(18) and B(53)) xor (A(19) and B(52)) xor (A(20) and B(51)) xor (A(21) and B(50)) xor (A(23) and B(49)) xor (A(23) and B(48)) xor (A(24) and B(47)) xor (A(25) and B(46)) xor (A(26) and B(45)) xor (A(27) and B(44)) xor (A(28) and B(43)) xor (A(29) and B(42)) xor (A(30) and B(41)) xor (A(31) and B(40)) xor (A(32) and B(39)) xor (A(33) and B(38)) xor (A(34) and B(37)) xor (A(35) and B(36)) xor (A(36) and B(35)) xor (A(37) and B(34)) xor (A(38) and B(33)) xor (A(39) and B(32)) xor (A(40) and B(31)) xor (A(41) and B(30)) xor (A(42) and B(29)) xor (A(43) and B(28)) xor (A(44) and B(27)) xor (A(45) and B(26)) xor (A(46) and B(25)) xor (A(47) and B(24)) xor (A(48) and B(23)) xor (A(49) and B(23)) xor (A(50) and B(21)) xor (A(51) and B(20)) xor (A(52) and B(19)) xor (A(53) and B(18)) xor (A(54) and B(17)) xor (A(55) and B(16)) xor (A(56) and B(15)) xor (A(57) and B(14)) xor (A(58) and B(13)) xor (A(59) and B(12)) xor (A(60) and B(11)) xor (A(61) and B(10)) xor (A(62) and B(9)) xor (A(63) and B(8)) xor (A(64) and B(7)) xor (A(65) and B(6)) xor (A(66) and B(5)) xor (A(67) and B(4)) xor (A(68) and B(3)) xor (A(69) and B(2)) xor (A(70) and B(1)) xor (A(71) and B(0)) xor (A(64) and B(127)) xor (A(65) and B(126)) xor (A(66) and B(125)) xor (A(67) and B(124)) xor (A(68) and B(123)) xor (A(69) and B(122)) xor (A(70) and B(121)) xor (A(71) and B(120)) xor (A(72) and B(119)) xor (A(73) and B(118)) xor (A(74) and B(117)) xor (A(75) and B(116)) xor (A(76) and B(115)) xor (A(77) and B(114)) xor (A(78) and B(113)) xor (A(79) and B(112)) xor (A(80) and B(111)) xor (A(81) and B(110)) xor (A(82) and B(109)) xor (A(83) and B(108)) xor (A(84) and B(107)) xor (A(85) and B(106)) xor (A(86) and B(105)) xor (A(87) and B(104)) xor (A(88) and B(103)) xor (A(89) and B(102)) xor (A(90) and B(101)) xor (A(91) and B(100)) xor (A(92) and B(99)) xor (A(93) and B(98)) xor (A(94) and B(97)) xor (A(95) and B(96)) xor (A(96) and B(95)) xor (A(97) and B(94)) xor (A(98) and B(93)) xor (A(99) and B(92)) xor (A(100) and B(91)) xor (A(101) and B(90)) xor (A(102) and B(89)) xor (A(103) and B(88)) xor (A(104) and B(87)) xor (A(105) and B(86)) xor (A(106) and B(85)) xor (A(107) and B(84)) xor (A(108) and B(83)) xor (A(109) and B(82)) xor (A(110) and B(81)) xor (A(111) and B(80)) xor (A(112) and B(79)) xor (A(113) and B(78)) xor (A(114) and B(77)) xor (A(115) and B(76)) xor (A(116) and B(75)) xor (A(117) and B(74)) xor (A(118) and B(73)) xor (A(119) and B(72)) xor (A(120) and B(71)) xor (A(121) and B(70)) xor (A(122) and B(69)) xor (A(123) and B(68)) xor (A(124) and B(67)) xor (A(125) and B(66)) xor (A(126) and B(65)) xor (A(69) and B(127)) xor (A(70) and B(126)) xor (A(71) and B(125)) xor (A(72) and B(124)) xor (A(73) and B(123)) xor (A(74) and B(122)) xor (A(75) and B(121)) xor (A(76) and B(120)) xor (A(77) and B(119)) xor (A(78) and B(118)) xor (A(79) and B(117)) xor (A(80) and B(116)) xor (A(81) and B(115)) xor (A(82) and B(114)) xor (A(83) and B(113)) xor (A(84) and B(112)) xor (A(85) and B(111)) xor (A(86) and B(110)) xor (A(87) and B(109)) xor (A(88) and B(108)) xor (A(89) and B(107)) xor (A(90) and B(106)) xor (A(91) and B(105)) xor (A(92) and B(104)) xor (A(93) and B(103)) xor (A(94) and B(102)) xor (A(95) and B(101)) xor (A(96) and B(100)) xor (A(97) and B(99)) xor (A(98) and B(98)) xor (A(99) and B(97)) xor (A(100) and B(96)) xor (A(101) and B(95)) xor (A(102) and B(94)) xor (A(103) and B(93)) xor (A(104) and B(92)) xor (A(105) and B(91)) xor (A(106) and B(90)) xor (A(107) and B(89)) xor (A(108) and B(88)) xor (A(109) and B(87)) xor (A(110) and B(86)) xor (A(111) and B(85)) xor (A(112) and B(84)) xor (A(113) and B(83)) xor (A(114) and B(82)) xor (A(115) and B(81)) xor (A(116) and B(80)) xor (A(117) and B(79)) xor (A(118) and B(78)) xor (A(119) and B(77)) xor (A(120) and B(76)) xor (A(121) and B(75)) xor (A(122) and B(74)) xor (A(123) and B(73)) xor (A(124) and B(72)) xor (A(125) and B(71)) xor (A(126) and B(70)) xor (A(70) and B(127)) xor (A(71) and B(126)) xor (A(72) and B(125)) xor (A(73) and B(124)) xor (A(74) and B(123)) xor (A(75) and B(122)) xor (A(76) and B(121)) xor (A(77) and B(120)) xor (A(78) and B(119)) xor (A(79) and B(118)) xor (A(80) and B(117)) xor (A(81) and B(116)) xor (A(82) and B(115)) xor (A(83) and B(114)) xor (A(84) and B(113)) xor (A(85) and B(112)) xor (A(86) and B(111)) xor (A(87) and B(110)) xor (A(88) and B(109)) xor (A(89) and B(108)) xor (A(90) and B(107)) xor (A(91) and B(106)) xor (A(92) and B(105)) xor (A(93) and B(104)) xor (A(94) and B(103)) xor (A(95) and B(102)) xor (A(96) and B(101)) xor (A(97) and B(100)) xor (A(98) and B(99)) xor (A(99) and B(98)) xor (A(100) and B(97)) xor (A(101) and B(96)) xor (A(102) and B(95)) xor (A(103) and B(94)) xor (A(104) and B(93)) xor (A(105) and B(92)) xor (A(106) and B(91)) xor (A(107) and B(90)) xor (A(108) and B(89)) xor (A(109) and B(88)) xor (A(110) and B(87)) xor (A(111) and B(86)) xor (A(112) and B(85)) xor (A(113) and B(84)) xor (A(114) and B(83)) xor (A(115) and B(82)) xor (A(116) and B(81)) xor (A(117) and B(80)) xor (A(118) and B(79)) xor (A(119) and B(78)) xor (A(120) and B(77)) xor (A(121) and B(76)) xor (A(122) and B(75)) xor (A(123) and B(74)) xor (A(124) and B(73)) xor (A(125) and B(72)) xor (A(126) and B(71)) xor (A(71) and B(127)) xor (A(72) and B(126)) xor (A(73) and B(125)) xor (A(74) and B(124)) xor (A(75) and B(123)) xor (A(76) and B(122)) xor (A(77) and B(121)) xor (A(78) and B(120)) xor (A(79) and B(119)) xor (A(80) and B(118)) xor (A(81) and B(117)) xor (A(82) and B(116)) xor (A(83) and B(115)) xor (A(84) and B(114)) xor (A(85) and B(113)) xor (A(86) and B(112)) xor (A(87) and B(111)) xor (A(88) and B(110)) xor (A(89) and B(109)) xor (A(90) and B(108)) xor (A(91) and B(107)) xor (A(92) and B(106)) xor (A(93) and B(105)) xor (A(94) and B(104)) xor (A(95) and B(103)) xor (A(96) and B(102)) xor (A(97) and B(101)) xor (A(98) and B(100)) xor (A(99) and B(99)) xor (A(100) and B(98)) xor (A(101) and B(97)) xor (A(102) and B(96)) xor (A(103) and B(95)) xor (A(104) and B(94)) xor (A(105) and B(93)) xor (A(106) and B(92)) xor (A(107) and B(91)) xor (A(108) and B(90)) xor (A(109) and B(89)) xor (A(110) and B(88)) xor (A(111) and B(87)) xor (A(112) and B(86)) xor (A(113) and B(85)) xor (A(114) and B(84)) xor (A(115) and B(83)) xor (A(116) and B(82)) xor (A(117) and B(81)) xor (A(118) and B(80)) xor (A(119) and B(79)) xor (A(120) and B(78)) xor (A(121) and B(77)) xor (A(122) and B(76)) xor (A(123) and B(75)) xor (A(124) and B(74)) xor (A(125) and B(73)) xor (A(126) and B(73));
    C(72)  <= (A(0) and B(72)) xor (A(1) and B(71)) xor (A(2) and B(70)) xor (A(3) and B(69)) xor (A(4) and B(68)) xor (A(5) and B(67)) xor (A(6) and B(66)) xor (A(7) and B(65)) xor (A(8) and B(64)) xor (A(9) and B(63)) xor (A(10) and B(62)) xor (A(11) and B(61)) xor (A(12) and B(60)) xor (A(13) and B(59)) xor (A(14) and B(58)) xor (A(15) and B(57)) xor (A(16) and B(56)) xor (A(17) and B(55)) xor (A(18) and B(54)) xor (A(19) and B(53)) xor (A(20) and B(52)) xor (A(21) and B(51)) xor (A(23) and B(50)) xor (A(23) and B(49)) xor (A(24) and B(48)) xor (A(25) and B(47)) xor (A(26) and B(46)) xor (A(27) and B(45)) xor (A(28) and B(44)) xor (A(29) and B(43)) xor (A(30) and B(42)) xor (A(31) and B(41)) xor (A(32) and B(40)) xor (A(33) and B(39)) xor (A(34) and B(38)) xor (A(35) and B(37)) xor (A(36) and B(36)) xor (A(37) and B(35)) xor (A(38) and B(34)) xor (A(39) and B(33)) xor (A(40) and B(32)) xor (A(41) and B(31)) xor (A(42) and B(30)) xor (A(43) and B(29)) xor (A(44) and B(28)) xor (A(45) and B(27)) xor (A(46) and B(26)) xor (A(47) and B(25)) xor (A(48) and B(24)) xor (A(49) and B(23)) xor (A(50) and B(23)) xor (A(51) and B(21)) xor (A(52) and B(20)) xor (A(53) and B(19)) xor (A(54) and B(18)) xor (A(55) and B(17)) xor (A(56) and B(16)) xor (A(57) and B(15)) xor (A(58) and B(14)) xor (A(59) and B(13)) xor (A(60) and B(12)) xor (A(61) and B(11)) xor (A(62) and B(10)) xor (A(63) and B(9)) xor (A(64) and B(8)) xor (A(65) and B(7)) xor (A(66) and B(6)) xor (A(67) and B(5)) xor (A(68) and B(4)) xor (A(69) and B(3)) xor (A(70) and B(2)) xor (A(71) and B(1)) xor (A(72) and B(0)) xor (A(65) and B(127)) xor (A(66) and B(126)) xor (A(67) and B(125)) xor (A(68) and B(124)) xor (A(69) and B(123)) xor (A(70) and B(122)) xor (A(71) and B(121)) xor (A(72) and B(120)) xor (A(73) and B(119)) xor (A(74) and B(118)) xor (A(75) and B(117)) xor (A(76) and B(116)) xor (A(77) and B(115)) xor (A(78) and B(114)) xor (A(79) and B(113)) xor (A(80) and B(112)) xor (A(81) and B(111)) xor (A(82) and B(110)) xor (A(83) and B(109)) xor (A(84) and B(108)) xor (A(85) and B(107)) xor (A(86) and B(106)) xor (A(87) and B(105)) xor (A(88) and B(104)) xor (A(89) and B(103)) xor (A(90) and B(102)) xor (A(91) and B(101)) xor (A(92) and B(100)) xor (A(93) and B(99)) xor (A(94) and B(98)) xor (A(95) and B(97)) xor (A(96) and B(96)) xor (A(97) and B(95)) xor (A(98) and B(94)) xor (A(99) and B(93)) xor (A(100) and B(92)) xor (A(101) and B(91)) xor (A(102) and B(90)) xor (A(103) and B(89)) xor (A(104) and B(88)) xor (A(105) and B(87)) xor (A(106) and B(86)) xor (A(107) and B(85)) xor (A(108) and B(84)) xor (A(109) and B(83)) xor (A(110) and B(82)) xor (A(111) and B(81)) xor (A(112) and B(80)) xor (A(113) and B(79)) xor (A(114) and B(78)) xor (A(115) and B(77)) xor (A(116) and B(76)) xor (A(117) and B(75)) xor (A(118) and B(74)) xor (A(119) and B(73)) xor (A(120) and B(72)) xor (A(121) and B(71)) xor (A(122) and B(70)) xor (A(123) and B(69)) xor (A(124) and B(68)) xor (A(125) and B(67)) xor (A(126) and B(66)) xor (A(70) and B(127)) xor (A(71) and B(126)) xor (A(72) and B(125)) xor (A(73) and B(124)) xor (A(74) and B(123)) xor (A(75) and B(122)) xor (A(76) and B(121)) xor (A(77) and B(120)) xor (A(78) and B(119)) xor (A(79) and B(118)) xor (A(80) and B(117)) xor (A(81) and B(116)) xor (A(82) and B(115)) xor (A(83) and B(114)) xor (A(84) and B(113)) xor (A(85) and B(112)) xor (A(86) and B(111)) xor (A(87) and B(110)) xor (A(88) and B(109)) xor (A(89) and B(108)) xor (A(90) and B(107)) xor (A(91) and B(106)) xor (A(92) and B(105)) xor (A(93) and B(104)) xor (A(94) and B(103)) xor (A(95) and B(102)) xor (A(96) and B(101)) xor (A(97) and B(100)) xor (A(98) and B(99)) xor (A(99) and B(98)) xor (A(100) and B(97)) xor (A(101) and B(96)) xor (A(102) and B(95)) xor (A(103) and B(94)) xor (A(104) and B(93)) xor (A(105) and B(92)) xor (A(106) and B(91)) xor (A(107) and B(90)) xor (A(108) and B(89)) xor (A(109) and B(88)) xor (A(110) and B(87)) xor (A(111) and B(86)) xor (A(112) and B(85)) xor (A(113) and B(84)) xor (A(114) and B(83)) xor (A(115) and B(82)) xor (A(116) and B(81)) xor (A(117) and B(80)) xor (A(118) and B(79)) xor (A(119) and B(78)) xor (A(120) and B(77)) xor (A(121) and B(76)) xor (A(122) and B(75)) xor (A(123) and B(74)) xor (A(124) and B(73)) xor (A(125) and B(72)) xor (A(126) and B(71)) xor (A(71) and B(127)) xor (A(72) and B(126)) xor (A(73) and B(125)) xor (A(74) and B(124)) xor (A(75) and B(123)) xor (A(76) and B(122)) xor (A(77) and B(121)) xor (A(78) and B(120)) xor (A(79) and B(119)) xor (A(80) and B(118)) xor (A(81) and B(117)) xor (A(82) and B(116)) xor (A(83) and B(115)) xor (A(84) and B(114)) xor (A(85) and B(113)) xor (A(86) and B(112)) xor (A(87) and B(111)) xor (A(88) and B(110)) xor (A(89) and B(109)) xor (A(90) and B(108)) xor (A(91) and B(107)) xor (A(92) and B(106)) xor (A(93) and B(105)) xor (A(94) and B(104)) xor (A(95) and B(103)) xor (A(96) and B(102)) xor (A(97) and B(101)) xor (A(98) and B(100)) xor (A(99) and B(99)) xor (A(100) and B(98)) xor (A(101) and B(97)) xor (A(102) and B(96)) xor (A(103) and B(95)) xor (A(104) and B(94)) xor (A(105) and B(93)) xor (A(106) and B(92)) xor (A(107) and B(91)) xor (A(108) and B(90)) xor (A(109) and B(89)) xor (A(110) and B(88)) xor (A(111) and B(87)) xor (A(112) and B(86)) xor (A(113) and B(85)) xor (A(114) and B(84)) xor (A(115) and B(83)) xor (A(116) and B(82)) xor (A(117) and B(81)) xor (A(118) and B(80)) xor (A(119) and B(79)) xor (A(120) and B(78)) xor (A(121) and B(77)) xor (A(122) and B(76)) xor (A(123) and B(75)) xor (A(124) and B(74)) xor (A(125) and B(73)) xor (A(126) and B(72)) xor (A(72) and B(127)) xor (A(73) and B(126)) xor (A(74) and B(125)) xor (A(75) and B(124)) xor (A(76) and B(123)) xor (A(77) and B(122)) xor (A(78) and B(121)) xor (A(79) and B(120)) xor (A(80) and B(119)) xor (A(81) and B(118)) xor (A(82) and B(117)) xor (A(83) and B(116)) xor (A(84) and B(115)) xor (A(85) and B(114)) xor (A(86) and B(113)) xor (A(87) and B(112)) xor (A(88) and B(111)) xor (A(89) and B(110)) xor (A(90) and B(109)) xor (A(91) and B(108)) xor (A(92) and B(107)) xor (A(93) and B(106)) xor (A(94) and B(105)) xor (A(95) and B(104)) xor (A(96) and B(103)) xor (A(97) and B(102)) xor (A(98) and B(101)) xor (A(99) and B(100)) xor (A(100) and B(99)) xor (A(101) and B(98)) xor (A(102) and B(97)) xor (A(103) and B(96)) xor (A(104) and B(95)) xor (A(105) and B(94)) xor (A(106) and B(93)) xor (A(107) and B(92)) xor (A(108) and B(91)) xor (A(109) and B(90)) xor (A(110) and B(89)) xor (A(111) and B(88)) xor (A(112) and B(87)) xor (A(113) and B(86)) xor (A(114) and B(85)) xor (A(115) and B(84)) xor (A(116) and B(83)) xor (A(117) and B(82)) xor (A(118) and B(81)) xor (A(119) and B(80)) xor (A(120) and B(79)) xor (A(121) and B(78)) xor (A(122) and B(77)) xor (A(123) and B(76)) xor (A(124) and B(75)) xor (A(125) and B(74)) xor (A(126) and B(74));
    C(73)  <= (A(0) and B(73)) xor (A(1) and B(72)) xor (A(2) and B(71)) xor (A(3) and B(70)) xor (A(4) and B(69)) xor (A(5) and B(68)) xor (A(6) and B(67)) xor (A(7) and B(66)) xor (A(8) and B(65)) xor (A(9) and B(64)) xor (A(10) and B(63)) xor (A(11) and B(62)) xor (A(12) and B(61)) xor (A(13) and B(60)) xor (A(14) and B(59)) xor (A(15) and B(58)) xor (A(16) and B(57)) xor (A(17) and B(56)) xor (A(18) and B(55)) xor (A(19) and B(54)) xor (A(20) and B(53)) xor (A(21) and B(52)) xor (A(23) and B(51)) xor (A(23) and B(50)) xor (A(24) and B(49)) xor (A(25) and B(48)) xor (A(26) and B(47)) xor (A(27) and B(46)) xor (A(28) and B(45)) xor (A(29) and B(44)) xor (A(30) and B(43)) xor (A(31) and B(42)) xor (A(32) and B(41)) xor (A(33) and B(40)) xor (A(34) and B(39)) xor (A(35) and B(38)) xor (A(36) and B(37)) xor (A(37) and B(36)) xor (A(38) and B(35)) xor (A(39) and B(34)) xor (A(40) and B(33)) xor (A(41) and B(32)) xor (A(42) and B(31)) xor (A(43) and B(30)) xor (A(44) and B(29)) xor (A(45) and B(28)) xor (A(46) and B(27)) xor (A(47) and B(26)) xor (A(48) and B(25)) xor (A(49) and B(24)) xor (A(50) and B(23)) xor (A(51) and B(23)) xor (A(52) and B(21)) xor (A(53) and B(20)) xor (A(54) and B(19)) xor (A(55) and B(18)) xor (A(56) and B(17)) xor (A(57) and B(16)) xor (A(58) and B(15)) xor (A(59) and B(14)) xor (A(60) and B(13)) xor (A(61) and B(12)) xor (A(62) and B(11)) xor (A(63) and B(10)) xor (A(64) and B(9)) xor (A(65) and B(8)) xor (A(66) and B(7)) xor (A(67) and B(6)) xor (A(68) and B(5)) xor (A(69) and B(4)) xor (A(70) and B(3)) xor (A(71) and B(2)) xor (A(72) and B(1)) xor (A(73) and B(0)) xor (A(66) and B(127)) xor (A(67) and B(126)) xor (A(68) and B(125)) xor (A(69) and B(124)) xor (A(70) and B(123)) xor (A(71) and B(122)) xor (A(72) and B(121)) xor (A(73) and B(120)) xor (A(74) and B(119)) xor (A(75) and B(118)) xor (A(76) and B(117)) xor (A(77) and B(116)) xor (A(78) and B(115)) xor (A(79) and B(114)) xor (A(80) and B(113)) xor (A(81) and B(112)) xor (A(82) and B(111)) xor (A(83) and B(110)) xor (A(84) and B(109)) xor (A(85) and B(108)) xor (A(86) and B(107)) xor (A(87) and B(106)) xor (A(88) and B(105)) xor (A(89) and B(104)) xor (A(90) and B(103)) xor (A(91) and B(102)) xor (A(92) and B(101)) xor (A(93) and B(100)) xor (A(94) and B(99)) xor (A(95) and B(98)) xor (A(96) and B(97)) xor (A(97) and B(96)) xor (A(98) and B(95)) xor (A(99) and B(94)) xor (A(100) and B(93)) xor (A(101) and B(92)) xor (A(102) and B(91)) xor (A(103) and B(90)) xor (A(104) and B(89)) xor (A(105) and B(88)) xor (A(106) and B(87)) xor (A(107) and B(86)) xor (A(108) and B(85)) xor (A(109) and B(84)) xor (A(110) and B(83)) xor (A(111) and B(82)) xor (A(112) and B(81)) xor (A(113) and B(80)) xor (A(114) and B(79)) xor (A(115) and B(78)) xor (A(116) and B(77)) xor (A(117) and B(76)) xor (A(118) and B(75)) xor (A(119) and B(74)) xor (A(120) and B(73)) xor (A(121) and B(72)) xor (A(122) and B(71)) xor (A(123) and B(70)) xor (A(124) and B(69)) xor (A(125) and B(68)) xor (A(126) and B(67)) xor (A(71) and B(127)) xor (A(72) and B(126)) xor (A(73) and B(125)) xor (A(74) and B(124)) xor (A(75) and B(123)) xor (A(76) and B(122)) xor (A(77) and B(121)) xor (A(78) and B(120)) xor (A(79) and B(119)) xor (A(80) and B(118)) xor (A(81) and B(117)) xor (A(82) and B(116)) xor (A(83) and B(115)) xor (A(84) and B(114)) xor (A(85) and B(113)) xor (A(86) and B(112)) xor (A(87) and B(111)) xor (A(88) and B(110)) xor (A(89) and B(109)) xor (A(90) and B(108)) xor (A(91) and B(107)) xor (A(92) and B(106)) xor (A(93) and B(105)) xor (A(94) and B(104)) xor (A(95) and B(103)) xor (A(96) and B(102)) xor (A(97) and B(101)) xor (A(98) and B(100)) xor (A(99) and B(99)) xor (A(100) and B(98)) xor (A(101) and B(97)) xor (A(102) and B(96)) xor (A(103) and B(95)) xor (A(104) and B(94)) xor (A(105) and B(93)) xor (A(106) and B(92)) xor (A(107) and B(91)) xor (A(108) and B(90)) xor (A(109) and B(89)) xor (A(110) and B(88)) xor (A(111) and B(87)) xor (A(112) and B(86)) xor (A(113) and B(85)) xor (A(114) and B(84)) xor (A(115) and B(83)) xor (A(116) and B(82)) xor (A(117) and B(81)) xor (A(118) and B(80)) xor (A(119) and B(79)) xor (A(120) and B(78)) xor (A(121) and B(77)) xor (A(122) and B(76)) xor (A(123) and B(75)) xor (A(124) and B(74)) xor (A(125) and B(73)) xor (A(126) and B(72)) xor (A(72) and B(127)) xor (A(73) and B(126)) xor (A(74) and B(125)) xor (A(75) and B(124)) xor (A(76) and B(123)) xor (A(77) and B(122)) xor (A(78) and B(121)) xor (A(79) and B(120)) xor (A(80) and B(119)) xor (A(81) and B(118)) xor (A(82) and B(117)) xor (A(83) and B(116)) xor (A(84) and B(115)) xor (A(85) and B(114)) xor (A(86) and B(113)) xor (A(87) and B(112)) xor (A(88) and B(111)) xor (A(89) and B(110)) xor (A(90) and B(109)) xor (A(91) and B(108)) xor (A(92) and B(107)) xor (A(93) and B(106)) xor (A(94) and B(105)) xor (A(95) and B(104)) xor (A(96) and B(103)) xor (A(97) and B(102)) xor (A(98) and B(101)) xor (A(99) and B(100)) xor (A(100) and B(99)) xor (A(101) and B(98)) xor (A(102) and B(97)) xor (A(103) and B(96)) xor (A(104) and B(95)) xor (A(105) and B(94)) xor (A(106) and B(93)) xor (A(107) and B(92)) xor (A(108) and B(91)) xor (A(109) and B(90)) xor (A(110) and B(89)) xor (A(111) and B(88)) xor (A(112) and B(87)) xor (A(113) and B(86)) xor (A(114) and B(85)) xor (A(115) and B(84)) xor (A(116) and B(83)) xor (A(117) and B(82)) xor (A(118) and B(81)) xor (A(119) and B(80)) xor (A(120) and B(79)) xor (A(121) and B(78)) xor (A(122) and B(77)) xor (A(123) and B(76)) xor (A(124) and B(75)) xor (A(125) and B(74)) xor (A(126) and B(73)) xor (A(73) and B(127)) xor (A(74) and B(126)) xor (A(75) and B(125)) xor (A(76) and B(124)) xor (A(77) and B(123)) xor (A(78) and B(122)) xor (A(79) and B(121)) xor (A(80) and B(120)) xor (A(81) and B(119)) xor (A(82) and B(118)) xor (A(83) and B(117)) xor (A(84) and B(116)) xor (A(85) and B(115)) xor (A(86) and B(114)) xor (A(87) and B(113)) xor (A(88) and B(112)) xor (A(89) and B(111)) xor (A(90) and B(110)) xor (A(91) and B(109)) xor (A(92) and B(108)) xor (A(93) and B(107)) xor (A(94) and B(106)) xor (A(95) and B(105)) xor (A(96) and B(104)) xor (A(97) and B(103)) xor (A(98) and B(102)) xor (A(99) and B(101)) xor (A(100) and B(100)) xor (A(101) and B(99)) xor (A(102) and B(98)) xor (A(103) and B(97)) xor (A(104) and B(96)) xor (A(105) and B(95)) xor (A(106) and B(94)) xor (A(107) and B(93)) xor (A(108) and B(92)) xor (A(109) and B(91)) xor (A(110) and B(90)) xor (A(111) and B(89)) xor (A(112) and B(88)) xor (A(113) and B(87)) xor (A(114) and B(86)) xor (A(115) and B(85)) xor (A(116) and B(84)) xor (A(117) and B(83)) xor (A(118) and B(82)) xor (A(119) and B(81)) xor (A(120) and B(80)) xor (A(121) and B(79)) xor (A(122) and B(78)) xor (A(123) and B(77)) xor (A(124) and B(76)) xor (A(125) and B(75)) xor (A(126) and B(75));
    C(74)  <= (A(0) and B(74)) xor (A(1) and B(73)) xor (A(2) and B(72)) xor (A(3) and B(71)) xor (A(4) and B(70)) xor (A(5) and B(69)) xor (A(6) and B(68)) xor (A(7) and B(67)) xor (A(8) and B(66)) xor (A(9) and B(65)) xor (A(10) and B(64)) xor (A(11) and B(63)) xor (A(12) and B(62)) xor (A(13) and B(61)) xor (A(14) and B(60)) xor (A(15) and B(59)) xor (A(16) and B(58)) xor (A(17) and B(57)) xor (A(18) and B(56)) xor (A(19) and B(55)) xor (A(20) and B(54)) xor (A(21) and B(53)) xor (A(23) and B(52)) xor (A(23) and B(51)) xor (A(24) and B(50)) xor (A(25) and B(49)) xor (A(26) and B(48)) xor (A(27) and B(47)) xor (A(28) and B(46)) xor (A(29) and B(45)) xor (A(30) and B(44)) xor (A(31) and B(43)) xor (A(32) and B(42)) xor (A(33) and B(41)) xor (A(34) and B(40)) xor (A(35) and B(39)) xor (A(36) and B(38)) xor (A(37) and B(37)) xor (A(38) and B(36)) xor (A(39) and B(35)) xor (A(40) and B(34)) xor (A(41) and B(33)) xor (A(42) and B(32)) xor (A(43) and B(31)) xor (A(44) and B(30)) xor (A(45) and B(29)) xor (A(46) and B(28)) xor (A(47) and B(27)) xor (A(48) and B(26)) xor (A(49) and B(25)) xor (A(50) and B(24)) xor (A(51) and B(23)) xor (A(52) and B(23)) xor (A(53) and B(21)) xor (A(54) and B(20)) xor (A(55) and B(19)) xor (A(56) and B(18)) xor (A(57) and B(17)) xor (A(58) and B(16)) xor (A(59) and B(15)) xor (A(60) and B(14)) xor (A(61) and B(13)) xor (A(62) and B(12)) xor (A(63) and B(11)) xor (A(64) and B(10)) xor (A(65) and B(9)) xor (A(66) and B(8)) xor (A(67) and B(7)) xor (A(68) and B(6)) xor (A(69) and B(5)) xor (A(70) and B(4)) xor (A(71) and B(3)) xor (A(72) and B(2)) xor (A(73) and B(1)) xor (A(74) and B(0)) xor (A(67) and B(127)) xor (A(68) and B(126)) xor (A(69) and B(125)) xor (A(70) and B(124)) xor (A(71) and B(123)) xor (A(72) and B(122)) xor (A(73) and B(121)) xor (A(74) and B(120)) xor (A(75) and B(119)) xor (A(76) and B(118)) xor (A(77) and B(117)) xor (A(78) and B(116)) xor (A(79) and B(115)) xor (A(80) and B(114)) xor (A(81) and B(113)) xor (A(82) and B(112)) xor (A(83) and B(111)) xor (A(84) and B(110)) xor (A(85) and B(109)) xor (A(86) and B(108)) xor (A(87) and B(107)) xor (A(88) and B(106)) xor (A(89) and B(105)) xor (A(90) and B(104)) xor (A(91) and B(103)) xor (A(92) and B(102)) xor (A(93) and B(101)) xor (A(94) and B(100)) xor (A(95) and B(99)) xor (A(96) and B(98)) xor (A(97) and B(97)) xor (A(98) and B(96)) xor (A(99) and B(95)) xor (A(100) and B(94)) xor (A(101) and B(93)) xor (A(102) and B(92)) xor (A(103) and B(91)) xor (A(104) and B(90)) xor (A(105) and B(89)) xor (A(106) and B(88)) xor (A(107) and B(87)) xor (A(108) and B(86)) xor (A(109) and B(85)) xor (A(110) and B(84)) xor (A(111) and B(83)) xor (A(112) and B(82)) xor (A(113) and B(81)) xor (A(114) and B(80)) xor (A(115) and B(79)) xor (A(116) and B(78)) xor (A(117) and B(77)) xor (A(118) and B(76)) xor (A(119) and B(75)) xor (A(120) and B(74)) xor (A(121) and B(73)) xor (A(122) and B(72)) xor (A(123) and B(71)) xor (A(124) and B(70)) xor (A(125) and B(69)) xor (A(126) and B(68)) xor (A(72) and B(127)) xor (A(73) and B(126)) xor (A(74) and B(125)) xor (A(75) and B(124)) xor (A(76) and B(123)) xor (A(77) and B(122)) xor (A(78) and B(121)) xor (A(79) and B(120)) xor (A(80) and B(119)) xor (A(81) and B(118)) xor (A(82) and B(117)) xor (A(83) and B(116)) xor (A(84) and B(115)) xor (A(85) and B(114)) xor (A(86) and B(113)) xor (A(87) and B(112)) xor (A(88) and B(111)) xor (A(89) and B(110)) xor (A(90) and B(109)) xor (A(91) and B(108)) xor (A(92) and B(107)) xor (A(93) and B(106)) xor (A(94) and B(105)) xor (A(95) and B(104)) xor (A(96) and B(103)) xor (A(97) and B(102)) xor (A(98) and B(101)) xor (A(99) and B(100)) xor (A(100) and B(99)) xor (A(101) and B(98)) xor (A(102) and B(97)) xor (A(103) and B(96)) xor (A(104) and B(95)) xor (A(105) and B(94)) xor (A(106) and B(93)) xor (A(107) and B(92)) xor (A(108) and B(91)) xor (A(109) and B(90)) xor (A(110) and B(89)) xor (A(111) and B(88)) xor (A(112) and B(87)) xor (A(113) and B(86)) xor (A(114) and B(85)) xor (A(115) and B(84)) xor (A(116) and B(83)) xor (A(117) and B(82)) xor (A(118) and B(81)) xor (A(119) and B(80)) xor (A(120) and B(79)) xor (A(121) and B(78)) xor (A(122) and B(77)) xor (A(123) and B(76)) xor (A(124) and B(75)) xor (A(125) and B(74)) xor (A(126) and B(73)) xor (A(73) and B(127)) xor (A(74) and B(126)) xor (A(75) and B(125)) xor (A(76) and B(124)) xor (A(77) and B(123)) xor (A(78) and B(122)) xor (A(79) and B(121)) xor (A(80) and B(120)) xor (A(81) and B(119)) xor (A(82) and B(118)) xor (A(83) and B(117)) xor (A(84) and B(116)) xor (A(85) and B(115)) xor (A(86) and B(114)) xor (A(87) and B(113)) xor (A(88) and B(112)) xor (A(89) and B(111)) xor (A(90) and B(110)) xor (A(91) and B(109)) xor (A(92) and B(108)) xor (A(93) and B(107)) xor (A(94) and B(106)) xor (A(95) and B(105)) xor (A(96) and B(104)) xor (A(97) and B(103)) xor (A(98) and B(102)) xor (A(99) and B(101)) xor (A(100) and B(100)) xor (A(101) and B(99)) xor (A(102) and B(98)) xor (A(103) and B(97)) xor (A(104) and B(96)) xor (A(105) and B(95)) xor (A(106) and B(94)) xor (A(107) and B(93)) xor (A(108) and B(92)) xor (A(109) and B(91)) xor (A(110) and B(90)) xor (A(111) and B(89)) xor (A(112) and B(88)) xor (A(113) and B(87)) xor (A(114) and B(86)) xor (A(115) and B(85)) xor (A(116) and B(84)) xor (A(117) and B(83)) xor (A(118) and B(82)) xor (A(119) and B(81)) xor (A(120) and B(80)) xor (A(121) and B(79)) xor (A(122) and B(78)) xor (A(123) and B(77)) xor (A(124) and B(76)) xor (A(125) and B(75)) xor (A(126) and B(74)) xor (A(74) and B(127)) xor (A(75) and B(126)) xor (A(76) and B(125)) xor (A(77) and B(124)) xor (A(78) and B(123)) xor (A(79) and B(122)) xor (A(80) and B(121)) xor (A(81) and B(120)) xor (A(82) and B(119)) xor (A(83) and B(118)) xor (A(84) and B(117)) xor (A(85) and B(116)) xor (A(86) and B(115)) xor (A(87) and B(114)) xor (A(88) and B(113)) xor (A(89) and B(112)) xor (A(90) and B(111)) xor (A(91) and B(110)) xor (A(92) and B(109)) xor (A(93) and B(108)) xor (A(94) and B(107)) xor (A(95) and B(106)) xor (A(96) and B(105)) xor (A(97) and B(104)) xor (A(98) and B(103)) xor (A(99) and B(102)) xor (A(100) and B(101)) xor (A(101) and B(100)) xor (A(102) and B(99)) xor (A(103) and B(98)) xor (A(104) and B(97)) xor (A(105) and B(96)) xor (A(106) and B(95)) xor (A(107) and B(94)) xor (A(108) and B(93)) xor (A(109) and B(92)) xor (A(110) and B(91)) xor (A(111) and B(90)) xor (A(112) and B(89)) xor (A(113) and B(88)) xor (A(114) and B(87)) xor (A(115) and B(86)) xor (A(116) and B(85)) xor (A(117) and B(84)) xor (A(118) and B(83)) xor (A(119) and B(82)) xor (A(120) and B(81)) xor (A(121) and B(80)) xor (A(122) and B(79)) xor (A(123) and B(78)) xor (A(124) and B(77)) xor (A(125) and B(76)) xor (A(126) and B(76));
    C(75)  <= (A(0) and B(75)) xor (A(1) and B(74)) xor (A(2) and B(73)) xor (A(3) and B(72)) xor (A(4) and B(71)) xor (A(5) and B(70)) xor (A(6) and B(69)) xor (A(7) and B(68)) xor (A(8) and B(67)) xor (A(9) and B(66)) xor (A(10) and B(65)) xor (A(11) and B(64)) xor (A(12) and B(63)) xor (A(13) and B(62)) xor (A(14) and B(61)) xor (A(15) and B(60)) xor (A(16) and B(59)) xor (A(17) and B(58)) xor (A(18) and B(57)) xor (A(19) and B(56)) xor (A(20) and B(55)) xor (A(21) and B(54)) xor (A(23) and B(53)) xor (A(23) and B(52)) xor (A(24) and B(51)) xor (A(25) and B(50)) xor (A(26) and B(49)) xor (A(27) and B(48)) xor (A(28) and B(47)) xor (A(29) and B(46)) xor (A(30) and B(45)) xor (A(31) and B(44)) xor (A(32) and B(43)) xor (A(33) and B(42)) xor (A(34) and B(41)) xor (A(35) and B(40)) xor (A(36) and B(39)) xor (A(37) and B(38)) xor (A(38) and B(37)) xor (A(39) and B(36)) xor (A(40) and B(35)) xor (A(41) and B(34)) xor (A(42) and B(33)) xor (A(43) and B(32)) xor (A(44) and B(31)) xor (A(45) and B(30)) xor (A(46) and B(29)) xor (A(47) and B(28)) xor (A(48) and B(27)) xor (A(49) and B(26)) xor (A(50) and B(25)) xor (A(51) and B(24)) xor (A(52) and B(23)) xor (A(53) and B(23)) xor (A(54) and B(21)) xor (A(55) and B(20)) xor (A(56) and B(19)) xor (A(57) and B(18)) xor (A(58) and B(17)) xor (A(59) and B(16)) xor (A(60) and B(15)) xor (A(61) and B(14)) xor (A(62) and B(13)) xor (A(63) and B(12)) xor (A(64) and B(11)) xor (A(65) and B(10)) xor (A(66) and B(9)) xor (A(67) and B(8)) xor (A(68) and B(7)) xor (A(69) and B(6)) xor (A(70) and B(5)) xor (A(71) and B(4)) xor (A(72) and B(3)) xor (A(73) and B(2)) xor (A(74) and B(1)) xor (A(75) and B(0)) xor (A(68) and B(127)) xor (A(69) and B(126)) xor (A(70) and B(125)) xor (A(71) and B(124)) xor (A(72) and B(123)) xor (A(73) and B(122)) xor (A(74) and B(121)) xor (A(75) and B(120)) xor (A(76) and B(119)) xor (A(77) and B(118)) xor (A(78) and B(117)) xor (A(79) and B(116)) xor (A(80) and B(115)) xor (A(81) and B(114)) xor (A(82) and B(113)) xor (A(83) and B(112)) xor (A(84) and B(111)) xor (A(85) and B(110)) xor (A(86) and B(109)) xor (A(87) and B(108)) xor (A(88) and B(107)) xor (A(89) and B(106)) xor (A(90) and B(105)) xor (A(91) and B(104)) xor (A(92) and B(103)) xor (A(93) and B(102)) xor (A(94) and B(101)) xor (A(95) and B(100)) xor (A(96) and B(99)) xor (A(97) and B(98)) xor (A(98) and B(97)) xor (A(99) and B(96)) xor (A(100) and B(95)) xor (A(101) and B(94)) xor (A(102) and B(93)) xor (A(103) and B(92)) xor (A(104) and B(91)) xor (A(105) and B(90)) xor (A(106) and B(89)) xor (A(107) and B(88)) xor (A(108) and B(87)) xor (A(109) and B(86)) xor (A(110) and B(85)) xor (A(111) and B(84)) xor (A(112) and B(83)) xor (A(113) and B(82)) xor (A(114) and B(81)) xor (A(115) and B(80)) xor (A(116) and B(79)) xor (A(117) and B(78)) xor (A(118) and B(77)) xor (A(119) and B(76)) xor (A(120) and B(75)) xor (A(121) and B(74)) xor (A(122) and B(73)) xor (A(123) and B(72)) xor (A(124) and B(71)) xor (A(125) and B(70)) xor (A(126) and B(69)) xor (A(73) and B(127)) xor (A(74) and B(126)) xor (A(75) and B(125)) xor (A(76) and B(124)) xor (A(77) and B(123)) xor (A(78) and B(122)) xor (A(79) and B(121)) xor (A(80) and B(120)) xor (A(81) and B(119)) xor (A(82) and B(118)) xor (A(83) and B(117)) xor (A(84) and B(116)) xor (A(85) and B(115)) xor (A(86) and B(114)) xor (A(87) and B(113)) xor (A(88) and B(112)) xor (A(89) and B(111)) xor (A(90) and B(110)) xor (A(91) and B(109)) xor (A(92) and B(108)) xor (A(93) and B(107)) xor (A(94) and B(106)) xor (A(95) and B(105)) xor (A(96) and B(104)) xor (A(97) and B(103)) xor (A(98) and B(102)) xor (A(99) and B(101)) xor (A(100) and B(100)) xor (A(101) and B(99)) xor (A(102) and B(98)) xor (A(103) and B(97)) xor (A(104) and B(96)) xor (A(105) and B(95)) xor (A(106) and B(94)) xor (A(107) and B(93)) xor (A(108) and B(92)) xor (A(109) and B(91)) xor (A(110) and B(90)) xor (A(111) and B(89)) xor (A(112) and B(88)) xor (A(113) and B(87)) xor (A(114) and B(86)) xor (A(115) and B(85)) xor (A(116) and B(84)) xor (A(117) and B(83)) xor (A(118) and B(82)) xor (A(119) and B(81)) xor (A(120) and B(80)) xor (A(121) and B(79)) xor (A(122) and B(78)) xor (A(123) and B(77)) xor (A(124) and B(76)) xor (A(125) and B(75)) xor (A(126) and B(74)) xor (A(74) and B(127)) xor (A(75) and B(126)) xor (A(76) and B(125)) xor (A(77) and B(124)) xor (A(78) and B(123)) xor (A(79) and B(122)) xor (A(80) and B(121)) xor (A(81) and B(120)) xor (A(82) and B(119)) xor (A(83) and B(118)) xor (A(84) and B(117)) xor (A(85) and B(116)) xor (A(86) and B(115)) xor (A(87) and B(114)) xor (A(88) and B(113)) xor (A(89) and B(112)) xor (A(90) and B(111)) xor (A(91) and B(110)) xor (A(92) and B(109)) xor (A(93) and B(108)) xor (A(94) and B(107)) xor (A(95) and B(106)) xor (A(96) and B(105)) xor (A(97) and B(104)) xor (A(98) and B(103)) xor (A(99) and B(102)) xor (A(100) and B(101)) xor (A(101) and B(100)) xor (A(102) and B(99)) xor (A(103) and B(98)) xor (A(104) and B(97)) xor (A(105) and B(96)) xor (A(106) and B(95)) xor (A(107) and B(94)) xor (A(108) and B(93)) xor (A(109) and B(92)) xor (A(110) and B(91)) xor (A(111) and B(90)) xor (A(112) and B(89)) xor (A(113) and B(88)) xor (A(114) and B(87)) xor (A(115) and B(86)) xor (A(116) and B(85)) xor (A(117) and B(84)) xor (A(118) and B(83)) xor (A(119) and B(82)) xor (A(120) and B(81)) xor (A(121) and B(80)) xor (A(122) and B(79)) xor (A(123) and B(78)) xor (A(124) and B(77)) xor (A(125) and B(76)) xor (A(126) and B(75)) xor (A(75) and B(127)) xor (A(76) and B(126)) xor (A(77) and B(125)) xor (A(78) and B(124)) xor (A(79) and B(123)) xor (A(80) and B(122)) xor (A(81) and B(121)) xor (A(82) and B(120)) xor (A(83) and B(119)) xor (A(84) and B(118)) xor (A(85) and B(117)) xor (A(86) and B(116)) xor (A(87) and B(115)) xor (A(88) and B(114)) xor (A(89) and B(113)) xor (A(90) and B(112)) xor (A(91) and B(111)) xor (A(92) and B(110)) xor (A(93) and B(109)) xor (A(94) and B(108)) xor (A(95) and B(107)) xor (A(96) and B(106)) xor (A(97) and B(105)) xor (A(98) and B(104)) xor (A(99) and B(103)) xor (A(100) and B(102)) xor (A(101) and B(101)) xor (A(102) and B(100)) xor (A(103) and B(99)) xor (A(104) and B(98)) xor (A(105) and B(97)) xor (A(106) and B(96)) xor (A(107) and B(95)) xor (A(108) and B(94)) xor (A(109) and B(93)) xor (A(110) and B(92)) xor (A(111) and B(91)) xor (A(112) and B(90)) xor (A(113) and B(89)) xor (A(114) and B(88)) xor (A(115) and B(87)) xor (A(116) and B(86)) xor (A(117) and B(85)) xor (A(118) and B(84)) xor (A(119) and B(83)) xor (A(120) and B(82)) xor (A(121) and B(81)) xor (A(122) and B(80)) xor (A(123) and B(79)) xor (A(124) and B(78)) xor (A(125) and B(77)) xor (A(126) and B(77));
    C(76)  <= (A(0) and B(76)) xor (A(1) and B(75)) xor (A(2) and B(74)) xor (A(3) and B(73)) xor (A(4) and B(72)) xor (A(5) and B(71)) xor (A(6) and B(70)) xor (A(7) and B(69)) xor (A(8) and B(68)) xor (A(9) and B(67)) xor (A(10) and B(66)) xor (A(11) and B(65)) xor (A(12) and B(64)) xor (A(13) and B(63)) xor (A(14) and B(62)) xor (A(15) and B(61)) xor (A(16) and B(60)) xor (A(17) and B(59)) xor (A(18) and B(58)) xor (A(19) and B(57)) xor (A(20) and B(56)) xor (A(21) and B(55)) xor (A(23) and B(54)) xor (A(23) and B(53)) xor (A(24) and B(52)) xor (A(25) and B(51)) xor (A(26) and B(50)) xor (A(27) and B(49)) xor (A(28) and B(48)) xor (A(29) and B(47)) xor (A(30) and B(46)) xor (A(31) and B(45)) xor (A(32) and B(44)) xor (A(33) and B(43)) xor (A(34) and B(42)) xor (A(35) and B(41)) xor (A(36) and B(40)) xor (A(37) and B(39)) xor (A(38) and B(38)) xor (A(39) and B(37)) xor (A(40) and B(36)) xor (A(41) and B(35)) xor (A(42) and B(34)) xor (A(43) and B(33)) xor (A(44) and B(32)) xor (A(45) and B(31)) xor (A(46) and B(30)) xor (A(47) and B(29)) xor (A(48) and B(28)) xor (A(49) and B(27)) xor (A(50) and B(26)) xor (A(51) and B(25)) xor (A(52) and B(24)) xor (A(53) and B(23)) xor (A(54) and B(23)) xor (A(55) and B(21)) xor (A(56) and B(20)) xor (A(57) and B(19)) xor (A(58) and B(18)) xor (A(59) and B(17)) xor (A(60) and B(16)) xor (A(61) and B(15)) xor (A(62) and B(14)) xor (A(63) and B(13)) xor (A(64) and B(12)) xor (A(65) and B(11)) xor (A(66) and B(10)) xor (A(67) and B(9)) xor (A(68) and B(8)) xor (A(69) and B(7)) xor (A(70) and B(6)) xor (A(71) and B(5)) xor (A(72) and B(4)) xor (A(73) and B(3)) xor (A(74) and B(2)) xor (A(75) and B(1)) xor (A(76) and B(0)) xor (A(69) and B(127)) xor (A(70) and B(126)) xor (A(71) and B(125)) xor (A(72) and B(124)) xor (A(73) and B(123)) xor (A(74) and B(122)) xor (A(75) and B(121)) xor (A(76) and B(120)) xor (A(77) and B(119)) xor (A(78) and B(118)) xor (A(79) and B(117)) xor (A(80) and B(116)) xor (A(81) and B(115)) xor (A(82) and B(114)) xor (A(83) and B(113)) xor (A(84) and B(112)) xor (A(85) and B(111)) xor (A(86) and B(110)) xor (A(87) and B(109)) xor (A(88) and B(108)) xor (A(89) and B(107)) xor (A(90) and B(106)) xor (A(91) and B(105)) xor (A(92) and B(104)) xor (A(93) and B(103)) xor (A(94) and B(102)) xor (A(95) and B(101)) xor (A(96) and B(100)) xor (A(97) and B(99)) xor (A(98) and B(98)) xor (A(99) and B(97)) xor (A(100) and B(96)) xor (A(101) and B(95)) xor (A(102) and B(94)) xor (A(103) and B(93)) xor (A(104) and B(92)) xor (A(105) and B(91)) xor (A(106) and B(90)) xor (A(107) and B(89)) xor (A(108) and B(88)) xor (A(109) and B(87)) xor (A(110) and B(86)) xor (A(111) and B(85)) xor (A(112) and B(84)) xor (A(113) and B(83)) xor (A(114) and B(82)) xor (A(115) and B(81)) xor (A(116) and B(80)) xor (A(117) and B(79)) xor (A(118) and B(78)) xor (A(119) and B(77)) xor (A(120) and B(76)) xor (A(121) and B(75)) xor (A(122) and B(74)) xor (A(123) and B(73)) xor (A(124) and B(72)) xor (A(125) and B(71)) xor (A(126) and B(70)) xor (A(74) and B(127)) xor (A(75) and B(126)) xor (A(76) and B(125)) xor (A(77) and B(124)) xor (A(78) and B(123)) xor (A(79) and B(122)) xor (A(80) and B(121)) xor (A(81) and B(120)) xor (A(82) and B(119)) xor (A(83) and B(118)) xor (A(84) and B(117)) xor (A(85) and B(116)) xor (A(86) and B(115)) xor (A(87) and B(114)) xor (A(88) and B(113)) xor (A(89) and B(112)) xor (A(90) and B(111)) xor (A(91) and B(110)) xor (A(92) and B(109)) xor (A(93) and B(108)) xor (A(94) and B(107)) xor (A(95) and B(106)) xor (A(96) and B(105)) xor (A(97) and B(104)) xor (A(98) and B(103)) xor (A(99) and B(102)) xor (A(100) and B(101)) xor (A(101) and B(100)) xor (A(102) and B(99)) xor (A(103) and B(98)) xor (A(104) and B(97)) xor (A(105) and B(96)) xor (A(106) and B(95)) xor (A(107) and B(94)) xor (A(108) and B(93)) xor (A(109) and B(92)) xor (A(110) and B(91)) xor (A(111) and B(90)) xor (A(112) and B(89)) xor (A(113) and B(88)) xor (A(114) and B(87)) xor (A(115) and B(86)) xor (A(116) and B(85)) xor (A(117) and B(84)) xor (A(118) and B(83)) xor (A(119) and B(82)) xor (A(120) and B(81)) xor (A(121) and B(80)) xor (A(122) and B(79)) xor (A(123) and B(78)) xor (A(124) and B(77)) xor (A(125) and B(76)) xor (A(126) and B(75)) xor (A(75) and B(127)) xor (A(76) and B(126)) xor (A(77) and B(125)) xor (A(78) and B(124)) xor (A(79) and B(123)) xor (A(80) and B(122)) xor (A(81) and B(121)) xor (A(82) and B(120)) xor (A(83) and B(119)) xor (A(84) and B(118)) xor (A(85) and B(117)) xor (A(86) and B(116)) xor (A(87) and B(115)) xor (A(88) and B(114)) xor (A(89) and B(113)) xor (A(90) and B(112)) xor (A(91) and B(111)) xor (A(92) and B(110)) xor (A(93) and B(109)) xor (A(94) and B(108)) xor (A(95) and B(107)) xor (A(96) and B(106)) xor (A(97) and B(105)) xor (A(98) and B(104)) xor (A(99) and B(103)) xor (A(100) and B(102)) xor (A(101) and B(101)) xor (A(102) and B(100)) xor (A(103) and B(99)) xor (A(104) and B(98)) xor (A(105) and B(97)) xor (A(106) and B(96)) xor (A(107) and B(95)) xor (A(108) and B(94)) xor (A(109) and B(93)) xor (A(110) and B(92)) xor (A(111) and B(91)) xor (A(112) and B(90)) xor (A(113) and B(89)) xor (A(114) and B(88)) xor (A(115) and B(87)) xor (A(116) and B(86)) xor (A(117) and B(85)) xor (A(118) and B(84)) xor (A(119) and B(83)) xor (A(120) and B(82)) xor (A(121) and B(81)) xor (A(122) and B(80)) xor (A(123) and B(79)) xor (A(124) and B(78)) xor (A(125) and B(77)) xor (A(126) and B(76)) xor (A(76) and B(127)) xor (A(77) and B(126)) xor (A(78) and B(125)) xor (A(79) and B(124)) xor (A(80) and B(123)) xor (A(81) and B(122)) xor (A(82) and B(121)) xor (A(83) and B(120)) xor (A(84) and B(119)) xor (A(85) and B(118)) xor (A(86) and B(117)) xor (A(87) and B(116)) xor (A(88) and B(115)) xor (A(89) and B(114)) xor (A(90) and B(113)) xor (A(91) and B(112)) xor (A(92) and B(111)) xor (A(93) and B(110)) xor (A(94) and B(109)) xor (A(95) and B(108)) xor (A(96) and B(107)) xor (A(97) and B(106)) xor (A(98) and B(105)) xor (A(99) and B(104)) xor (A(100) and B(103)) xor (A(101) and B(102)) xor (A(102) and B(101)) xor (A(103) and B(100)) xor (A(104) and B(99)) xor (A(105) and B(98)) xor (A(106) and B(97)) xor (A(107) and B(96)) xor (A(108) and B(95)) xor (A(109) and B(94)) xor (A(110) and B(93)) xor (A(111) and B(92)) xor (A(112) and B(91)) xor (A(113) and B(90)) xor (A(114) and B(89)) xor (A(115) and B(88)) xor (A(116) and B(87)) xor (A(117) and B(86)) xor (A(118) and B(85)) xor (A(119) and B(84)) xor (A(120) and B(83)) xor (A(121) and B(82)) xor (A(122) and B(81)) xor (A(123) and B(80)) xor (A(124) and B(79)) xor (A(125) and B(78)) xor (A(126) and B(78));
    C(77)  <= (A(0) and B(77)) xor (A(1) and B(76)) xor (A(2) and B(75)) xor (A(3) and B(74)) xor (A(4) and B(73)) xor (A(5) and B(72)) xor (A(6) and B(71)) xor (A(7) and B(70)) xor (A(8) and B(69)) xor (A(9) and B(68)) xor (A(10) and B(67)) xor (A(11) and B(66)) xor (A(12) and B(65)) xor (A(13) and B(64)) xor (A(14) and B(63)) xor (A(15) and B(62)) xor (A(16) and B(61)) xor (A(17) and B(60)) xor (A(18) and B(59)) xor (A(19) and B(58)) xor (A(20) and B(57)) xor (A(21) and B(56)) xor (A(23) and B(55)) xor (A(23) and B(54)) xor (A(24) and B(53)) xor (A(25) and B(52)) xor (A(26) and B(51)) xor (A(27) and B(50)) xor (A(28) and B(49)) xor (A(29) and B(48)) xor (A(30) and B(47)) xor (A(31) and B(46)) xor (A(32) and B(45)) xor (A(33) and B(44)) xor (A(34) and B(43)) xor (A(35) and B(42)) xor (A(36) and B(41)) xor (A(37) and B(40)) xor (A(38) and B(39)) xor (A(39) and B(38)) xor (A(40) and B(37)) xor (A(41) and B(36)) xor (A(42) and B(35)) xor (A(43) and B(34)) xor (A(44) and B(33)) xor (A(45) and B(32)) xor (A(46) and B(31)) xor (A(47) and B(30)) xor (A(48) and B(29)) xor (A(49) and B(28)) xor (A(50) and B(27)) xor (A(51) and B(26)) xor (A(52) and B(25)) xor (A(53) and B(24)) xor (A(54) and B(23)) xor (A(55) and B(23)) xor (A(56) and B(21)) xor (A(57) and B(20)) xor (A(58) and B(19)) xor (A(59) and B(18)) xor (A(60) and B(17)) xor (A(61) and B(16)) xor (A(62) and B(15)) xor (A(63) and B(14)) xor (A(64) and B(13)) xor (A(65) and B(12)) xor (A(66) and B(11)) xor (A(67) and B(10)) xor (A(68) and B(9)) xor (A(69) and B(8)) xor (A(70) and B(7)) xor (A(71) and B(6)) xor (A(72) and B(5)) xor (A(73) and B(4)) xor (A(74) and B(3)) xor (A(75) and B(2)) xor (A(76) and B(1)) xor (A(77) and B(0)) xor (A(70) and B(127)) xor (A(71) and B(126)) xor (A(72) and B(125)) xor (A(73) and B(124)) xor (A(74) and B(123)) xor (A(75) and B(122)) xor (A(76) and B(121)) xor (A(77) and B(120)) xor (A(78) and B(119)) xor (A(79) and B(118)) xor (A(80) and B(117)) xor (A(81) and B(116)) xor (A(82) and B(115)) xor (A(83) and B(114)) xor (A(84) and B(113)) xor (A(85) and B(112)) xor (A(86) and B(111)) xor (A(87) and B(110)) xor (A(88) and B(109)) xor (A(89) and B(108)) xor (A(90) and B(107)) xor (A(91) and B(106)) xor (A(92) and B(105)) xor (A(93) and B(104)) xor (A(94) and B(103)) xor (A(95) and B(102)) xor (A(96) and B(101)) xor (A(97) and B(100)) xor (A(98) and B(99)) xor (A(99) and B(98)) xor (A(100) and B(97)) xor (A(101) and B(96)) xor (A(102) and B(95)) xor (A(103) and B(94)) xor (A(104) and B(93)) xor (A(105) and B(92)) xor (A(106) and B(91)) xor (A(107) and B(90)) xor (A(108) and B(89)) xor (A(109) and B(88)) xor (A(110) and B(87)) xor (A(111) and B(86)) xor (A(112) and B(85)) xor (A(113) and B(84)) xor (A(114) and B(83)) xor (A(115) and B(82)) xor (A(116) and B(81)) xor (A(117) and B(80)) xor (A(118) and B(79)) xor (A(119) and B(78)) xor (A(120) and B(77)) xor (A(121) and B(76)) xor (A(122) and B(75)) xor (A(123) and B(74)) xor (A(124) and B(73)) xor (A(125) and B(72)) xor (A(126) and B(71)) xor (A(75) and B(127)) xor (A(76) and B(126)) xor (A(77) and B(125)) xor (A(78) and B(124)) xor (A(79) and B(123)) xor (A(80) and B(122)) xor (A(81) and B(121)) xor (A(82) and B(120)) xor (A(83) and B(119)) xor (A(84) and B(118)) xor (A(85) and B(117)) xor (A(86) and B(116)) xor (A(87) and B(115)) xor (A(88) and B(114)) xor (A(89) and B(113)) xor (A(90) and B(112)) xor (A(91) and B(111)) xor (A(92) and B(110)) xor (A(93) and B(109)) xor (A(94) and B(108)) xor (A(95) and B(107)) xor (A(96) and B(106)) xor (A(97) and B(105)) xor (A(98) and B(104)) xor (A(99) and B(103)) xor (A(100) and B(102)) xor (A(101) and B(101)) xor (A(102) and B(100)) xor (A(103) and B(99)) xor (A(104) and B(98)) xor (A(105) and B(97)) xor (A(106) and B(96)) xor (A(107) and B(95)) xor (A(108) and B(94)) xor (A(109) and B(93)) xor (A(110) and B(92)) xor (A(111) and B(91)) xor (A(112) and B(90)) xor (A(113) and B(89)) xor (A(114) and B(88)) xor (A(115) and B(87)) xor (A(116) and B(86)) xor (A(117) and B(85)) xor (A(118) and B(84)) xor (A(119) and B(83)) xor (A(120) and B(82)) xor (A(121) and B(81)) xor (A(122) and B(80)) xor (A(123) and B(79)) xor (A(124) and B(78)) xor (A(125) and B(77)) xor (A(126) and B(76)) xor (A(76) and B(127)) xor (A(77) and B(126)) xor (A(78) and B(125)) xor (A(79) and B(124)) xor (A(80) and B(123)) xor (A(81) and B(122)) xor (A(82) and B(121)) xor (A(83) and B(120)) xor (A(84) and B(119)) xor (A(85) and B(118)) xor (A(86) and B(117)) xor (A(87) and B(116)) xor (A(88) and B(115)) xor (A(89) and B(114)) xor (A(90) and B(113)) xor (A(91) and B(112)) xor (A(92) and B(111)) xor (A(93) and B(110)) xor (A(94) and B(109)) xor (A(95) and B(108)) xor (A(96) and B(107)) xor (A(97) and B(106)) xor (A(98) and B(105)) xor (A(99) and B(104)) xor (A(100) and B(103)) xor (A(101) and B(102)) xor (A(102) and B(101)) xor (A(103) and B(100)) xor (A(104) and B(99)) xor (A(105) and B(98)) xor (A(106) and B(97)) xor (A(107) and B(96)) xor (A(108) and B(95)) xor (A(109) and B(94)) xor (A(110) and B(93)) xor (A(111) and B(92)) xor (A(112) and B(91)) xor (A(113) and B(90)) xor (A(114) and B(89)) xor (A(115) and B(88)) xor (A(116) and B(87)) xor (A(117) and B(86)) xor (A(118) and B(85)) xor (A(119) and B(84)) xor (A(120) and B(83)) xor (A(121) and B(82)) xor (A(122) and B(81)) xor (A(123) and B(80)) xor (A(124) and B(79)) xor (A(125) and B(78)) xor (A(126) and B(77)) xor (A(77) and B(127)) xor (A(78) and B(126)) xor (A(79) and B(125)) xor (A(80) and B(124)) xor (A(81) and B(123)) xor (A(82) and B(122)) xor (A(83) and B(121)) xor (A(84) and B(120)) xor (A(85) and B(119)) xor (A(86) and B(118)) xor (A(87) and B(117)) xor (A(88) and B(116)) xor (A(89) and B(115)) xor (A(90) and B(114)) xor (A(91) and B(113)) xor (A(92) and B(112)) xor (A(93) and B(111)) xor (A(94) and B(110)) xor (A(95) and B(109)) xor (A(96) and B(108)) xor (A(97) and B(107)) xor (A(98) and B(106)) xor (A(99) and B(105)) xor (A(100) and B(104)) xor (A(101) and B(103)) xor (A(102) and B(102)) xor (A(103) and B(101)) xor (A(104) and B(100)) xor (A(105) and B(99)) xor (A(106) and B(98)) xor (A(107) and B(97)) xor (A(108) and B(96)) xor (A(109) and B(95)) xor (A(110) and B(94)) xor (A(111) and B(93)) xor (A(112) and B(92)) xor (A(113) and B(91)) xor (A(114) and B(90)) xor (A(115) and B(89)) xor (A(116) and B(88)) xor (A(117) and B(87)) xor (A(118) and B(86)) xor (A(119) and B(85)) xor (A(120) and B(84)) xor (A(121) and B(83)) xor (A(122) and B(82)) xor (A(123) and B(81)) xor (A(124) and B(80)) xor (A(125) and B(79)) xor (A(126) and B(79));
    C(78)  <= (A(0) and B(78)) xor (A(1) and B(77)) xor (A(2) and B(76)) xor (A(3) and B(75)) xor (A(4) and B(74)) xor (A(5) and B(73)) xor (A(6) and B(72)) xor (A(7) and B(71)) xor (A(8) and B(70)) xor (A(9) and B(69)) xor (A(10) and B(68)) xor (A(11) and B(67)) xor (A(12) and B(66)) xor (A(13) and B(65)) xor (A(14) and B(64)) xor (A(15) and B(63)) xor (A(16) and B(62)) xor (A(17) and B(61)) xor (A(18) and B(60)) xor (A(19) and B(59)) xor (A(20) and B(58)) xor (A(21) and B(57)) xor (A(23) and B(56)) xor (A(23) and B(55)) xor (A(24) and B(54)) xor (A(25) and B(53)) xor (A(26) and B(52)) xor (A(27) and B(51)) xor (A(28) and B(50)) xor (A(29) and B(49)) xor (A(30) and B(48)) xor (A(31) and B(47)) xor (A(32) and B(46)) xor (A(33) and B(45)) xor (A(34) and B(44)) xor (A(35) and B(43)) xor (A(36) and B(42)) xor (A(37) and B(41)) xor (A(38) and B(40)) xor (A(39) and B(39)) xor (A(40) and B(38)) xor (A(41) and B(37)) xor (A(42) and B(36)) xor (A(43) and B(35)) xor (A(44) and B(34)) xor (A(45) and B(33)) xor (A(46) and B(32)) xor (A(47) and B(31)) xor (A(48) and B(30)) xor (A(49) and B(29)) xor (A(50) and B(28)) xor (A(51) and B(27)) xor (A(52) and B(26)) xor (A(53) and B(25)) xor (A(54) and B(24)) xor (A(55) and B(23)) xor (A(56) and B(23)) xor (A(57) and B(21)) xor (A(58) and B(20)) xor (A(59) and B(19)) xor (A(60) and B(18)) xor (A(61) and B(17)) xor (A(62) and B(16)) xor (A(63) and B(15)) xor (A(64) and B(14)) xor (A(65) and B(13)) xor (A(66) and B(12)) xor (A(67) and B(11)) xor (A(68) and B(10)) xor (A(69) and B(9)) xor (A(70) and B(8)) xor (A(71) and B(7)) xor (A(72) and B(6)) xor (A(73) and B(5)) xor (A(74) and B(4)) xor (A(75) and B(3)) xor (A(76) and B(2)) xor (A(77) and B(1)) xor (A(78) and B(0)) xor (A(71) and B(127)) xor (A(72) and B(126)) xor (A(73) and B(125)) xor (A(74) and B(124)) xor (A(75) and B(123)) xor (A(76) and B(122)) xor (A(77) and B(121)) xor (A(78) and B(120)) xor (A(79) and B(119)) xor (A(80) and B(118)) xor (A(81) and B(117)) xor (A(82) and B(116)) xor (A(83) and B(115)) xor (A(84) and B(114)) xor (A(85) and B(113)) xor (A(86) and B(112)) xor (A(87) and B(111)) xor (A(88) and B(110)) xor (A(89) and B(109)) xor (A(90) and B(108)) xor (A(91) and B(107)) xor (A(92) and B(106)) xor (A(93) and B(105)) xor (A(94) and B(104)) xor (A(95) and B(103)) xor (A(96) and B(102)) xor (A(97) and B(101)) xor (A(98) and B(100)) xor (A(99) and B(99)) xor (A(100) and B(98)) xor (A(101) and B(97)) xor (A(102) and B(96)) xor (A(103) and B(95)) xor (A(104) and B(94)) xor (A(105) and B(93)) xor (A(106) and B(92)) xor (A(107) and B(91)) xor (A(108) and B(90)) xor (A(109) and B(89)) xor (A(110) and B(88)) xor (A(111) and B(87)) xor (A(112) and B(86)) xor (A(113) and B(85)) xor (A(114) and B(84)) xor (A(115) and B(83)) xor (A(116) and B(82)) xor (A(117) and B(81)) xor (A(118) and B(80)) xor (A(119) and B(79)) xor (A(120) and B(78)) xor (A(121) and B(77)) xor (A(122) and B(76)) xor (A(123) and B(75)) xor (A(124) and B(74)) xor (A(125) and B(73)) xor (A(126) and B(72)) xor (A(76) and B(127)) xor (A(77) and B(126)) xor (A(78) and B(125)) xor (A(79) and B(124)) xor (A(80) and B(123)) xor (A(81) and B(122)) xor (A(82) and B(121)) xor (A(83) and B(120)) xor (A(84) and B(119)) xor (A(85) and B(118)) xor (A(86) and B(117)) xor (A(87) and B(116)) xor (A(88) and B(115)) xor (A(89) and B(114)) xor (A(90) and B(113)) xor (A(91) and B(112)) xor (A(92) and B(111)) xor (A(93) and B(110)) xor (A(94) and B(109)) xor (A(95) and B(108)) xor (A(96) and B(107)) xor (A(97) and B(106)) xor (A(98) and B(105)) xor (A(99) and B(104)) xor (A(100) and B(103)) xor (A(101) and B(102)) xor (A(102) and B(101)) xor (A(103) and B(100)) xor (A(104) and B(99)) xor (A(105) and B(98)) xor (A(106) and B(97)) xor (A(107) and B(96)) xor (A(108) and B(95)) xor (A(109) and B(94)) xor (A(110) and B(93)) xor (A(111) and B(92)) xor (A(112) and B(91)) xor (A(113) and B(90)) xor (A(114) and B(89)) xor (A(115) and B(88)) xor (A(116) and B(87)) xor (A(117) and B(86)) xor (A(118) and B(85)) xor (A(119) and B(84)) xor (A(120) and B(83)) xor (A(121) and B(82)) xor (A(122) and B(81)) xor (A(123) and B(80)) xor (A(124) and B(79)) xor (A(125) and B(78)) xor (A(126) and B(77)) xor (A(77) and B(127)) xor (A(78) and B(126)) xor (A(79) and B(125)) xor (A(80) and B(124)) xor (A(81) and B(123)) xor (A(82) and B(122)) xor (A(83) and B(121)) xor (A(84) and B(120)) xor (A(85) and B(119)) xor (A(86) and B(118)) xor (A(87) and B(117)) xor (A(88) and B(116)) xor (A(89) and B(115)) xor (A(90) and B(114)) xor (A(91) and B(113)) xor (A(92) and B(112)) xor (A(93) and B(111)) xor (A(94) and B(110)) xor (A(95) and B(109)) xor (A(96) and B(108)) xor (A(97) and B(107)) xor (A(98) and B(106)) xor (A(99) and B(105)) xor (A(100) and B(104)) xor (A(101) and B(103)) xor (A(102) and B(102)) xor (A(103) and B(101)) xor (A(104) and B(100)) xor (A(105) and B(99)) xor (A(106) and B(98)) xor (A(107) and B(97)) xor (A(108) and B(96)) xor (A(109) and B(95)) xor (A(110) and B(94)) xor (A(111) and B(93)) xor (A(112) and B(92)) xor (A(113) and B(91)) xor (A(114) and B(90)) xor (A(115) and B(89)) xor (A(116) and B(88)) xor (A(117) and B(87)) xor (A(118) and B(86)) xor (A(119) and B(85)) xor (A(120) and B(84)) xor (A(121) and B(83)) xor (A(122) and B(82)) xor (A(123) and B(81)) xor (A(124) and B(80)) xor (A(125) and B(79)) xor (A(126) and B(78)) xor (A(78) and B(127)) xor (A(79) and B(126)) xor (A(80) and B(125)) xor (A(81) and B(124)) xor (A(82) and B(123)) xor (A(83) and B(122)) xor (A(84) and B(121)) xor (A(85) and B(120)) xor (A(86) and B(119)) xor (A(87) and B(118)) xor (A(88) and B(117)) xor (A(89) and B(116)) xor (A(90) and B(115)) xor (A(91) and B(114)) xor (A(92) and B(113)) xor (A(93) and B(112)) xor (A(94) and B(111)) xor (A(95) and B(110)) xor (A(96) and B(109)) xor (A(97) and B(108)) xor (A(98) and B(107)) xor (A(99) and B(106)) xor (A(100) and B(105)) xor (A(101) and B(104)) xor (A(102) and B(103)) xor (A(103) and B(102)) xor (A(104) and B(101)) xor (A(105) and B(100)) xor (A(106) and B(99)) xor (A(107) and B(98)) xor (A(108) and B(97)) xor (A(109) and B(96)) xor (A(110) and B(95)) xor (A(111) and B(94)) xor (A(112) and B(93)) xor (A(113) and B(92)) xor (A(114) and B(91)) xor (A(115) and B(90)) xor (A(116) and B(89)) xor (A(117) and B(88)) xor (A(118) and B(87)) xor (A(119) and B(86)) xor (A(120) and B(85)) xor (A(121) and B(84)) xor (A(122) and B(83)) xor (A(123) and B(82)) xor (A(124) and B(81)) xor (A(125) and B(80)) xor (A(126) and B(80));
    C(79)  <= (A(0) and B(79)) xor (A(1) and B(78)) xor (A(2) and B(77)) xor (A(3) and B(76)) xor (A(4) and B(75)) xor (A(5) and B(74)) xor (A(6) and B(73)) xor (A(7) and B(72)) xor (A(8) and B(71)) xor (A(9) and B(70)) xor (A(10) and B(69)) xor (A(11) and B(68)) xor (A(12) and B(67)) xor (A(13) and B(66)) xor (A(14) and B(65)) xor (A(15) and B(64)) xor (A(16) and B(63)) xor (A(17) and B(62)) xor (A(18) and B(61)) xor (A(19) and B(60)) xor (A(20) and B(59)) xor (A(21) and B(58)) xor (A(23) and B(57)) xor (A(23) and B(56)) xor (A(24) and B(55)) xor (A(25) and B(54)) xor (A(26) and B(53)) xor (A(27) and B(52)) xor (A(28) and B(51)) xor (A(29) and B(50)) xor (A(30) and B(49)) xor (A(31) and B(48)) xor (A(32) and B(47)) xor (A(33) and B(46)) xor (A(34) and B(45)) xor (A(35) and B(44)) xor (A(36) and B(43)) xor (A(37) and B(42)) xor (A(38) and B(41)) xor (A(39) and B(40)) xor (A(40) and B(39)) xor (A(41) and B(38)) xor (A(42) and B(37)) xor (A(43) and B(36)) xor (A(44) and B(35)) xor (A(45) and B(34)) xor (A(46) and B(33)) xor (A(47) and B(32)) xor (A(48) and B(31)) xor (A(49) and B(30)) xor (A(50) and B(29)) xor (A(51) and B(28)) xor (A(52) and B(27)) xor (A(53) and B(26)) xor (A(54) and B(25)) xor (A(55) and B(24)) xor (A(56) and B(23)) xor (A(57) and B(23)) xor (A(58) and B(21)) xor (A(59) and B(20)) xor (A(60) and B(19)) xor (A(61) and B(18)) xor (A(62) and B(17)) xor (A(63) and B(16)) xor (A(64) and B(15)) xor (A(65) and B(14)) xor (A(66) and B(13)) xor (A(67) and B(12)) xor (A(68) and B(11)) xor (A(69) and B(10)) xor (A(70) and B(9)) xor (A(71) and B(8)) xor (A(72) and B(7)) xor (A(73) and B(6)) xor (A(74) and B(5)) xor (A(75) and B(4)) xor (A(76) and B(3)) xor (A(77) and B(2)) xor (A(78) and B(1)) xor (A(79) and B(0)) xor (A(72) and B(127)) xor (A(73) and B(126)) xor (A(74) and B(125)) xor (A(75) and B(124)) xor (A(76) and B(123)) xor (A(77) and B(122)) xor (A(78) and B(121)) xor (A(79) and B(120)) xor (A(80) and B(119)) xor (A(81) and B(118)) xor (A(82) and B(117)) xor (A(83) and B(116)) xor (A(84) and B(115)) xor (A(85) and B(114)) xor (A(86) and B(113)) xor (A(87) and B(112)) xor (A(88) and B(111)) xor (A(89) and B(110)) xor (A(90) and B(109)) xor (A(91) and B(108)) xor (A(92) and B(107)) xor (A(93) and B(106)) xor (A(94) and B(105)) xor (A(95) and B(104)) xor (A(96) and B(103)) xor (A(97) and B(102)) xor (A(98) and B(101)) xor (A(99) and B(100)) xor (A(100) and B(99)) xor (A(101) and B(98)) xor (A(102) and B(97)) xor (A(103) and B(96)) xor (A(104) and B(95)) xor (A(105) and B(94)) xor (A(106) and B(93)) xor (A(107) and B(92)) xor (A(108) and B(91)) xor (A(109) and B(90)) xor (A(110) and B(89)) xor (A(111) and B(88)) xor (A(112) and B(87)) xor (A(113) and B(86)) xor (A(114) and B(85)) xor (A(115) and B(84)) xor (A(116) and B(83)) xor (A(117) and B(82)) xor (A(118) and B(81)) xor (A(119) and B(80)) xor (A(120) and B(79)) xor (A(121) and B(78)) xor (A(122) and B(77)) xor (A(123) and B(76)) xor (A(124) and B(75)) xor (A(125) and B(74)) xor (A(126) and B(73)) xor (A(77) and B(127)) xor (A(78) and B(126)) xor (A(79) and B(125)) xor (A(80) and B(124)) xor (A(81) and B(123)) xor (A(82) and B(122)) xor (A(83) and B(121)) xor (A(84) and B(120)) xor (A(85) and B(119)) xor (A(86) and B(118)) xor (A(87) and B(117)) xor (A(88) and B(116)) xor (A(89) and B(115)) xor (A(90) and B(114)) xor (A(91) and B(113)) xor (A(92) and B(112)) xor (A(93) and B(111)) xor (A(94) and B(110)) xor (A(95) and B(109)) xor (A(96) and B(108)) xor (A(97) and B(107)) xor (A(98) and B(106)) xor (A(99) and B(105)) xor (A(100) and B(104)) xor (A(101) and B(103)) xor (A(102) and B(102)) xor (A(103) and B(101)) xor (A(104) and B(100)) xor (A(105) and B(99)) xor (A(106) and B(98)) xor (A(107) and B(97)) xor (A(108) and B(96)) xor (A(109) and B(95)) xor (A(110) and B(94)) xor (A(111) and B(93)) xor (A(112) and B(92)) xor (A(113) and B(91)) xor (A(114) and B(90)) xor (A(115) and B(89)) xor (A(116) and B(88)) xor (A(117) and B(87)) xor (A(118) and B(86)) xor (A(119) and B(85)) xor (A(120) and B(84)) xor (A(121) and B(83)) xor (A(122) and B(82)) xor (A(123) and B(81)) xor (A(124) and B(80)) xor (A(125) and B(79)) xor (A(126) and B(78)) xor (A(78) and B(127)) xor (A(79) and B(126)) xor (A(80) and B(125)) xor (A(81) and B(124)) xor (A(82) and B(123)) xor (A(83) and B(122)) xor (A(84) and B(121)) xor (A(85) and B(120)) xor (A(86) and B(119)) xor (A(87) and B(118)) xor (A(88) and B(117)) xor (A(89) and B(116)) xor (A(90) and B(115)) xor (A(91) and B(114)) xor (A(92) and B(113)) xor (A(93) and B(112)) xor (A(94) and B(111)) xor (A(95) and B(110)) xor (A(96) and B(109)) xor (A(97) and B(108)) xor (A(98) and B(107)) xor (A(99) and B(106)) xor (A(100) and B(105)) xor (A(101) and B(104)) xor (A(102) and B(103)) xor (A(103) and B(102)) xor (A(104) and B(101)) xor (A(105) and B(100)) xor (A(106) and B(99)) xor (A(107) and B(98)) xor (A(108) and B(97)) xor (A(109) and B(96)) xor (A(110) and B(95)) xor (A(111) and B(94)) xor (A(112) and B(93)) xor (A(113) and B(92)) xor (A(114) and B(91)) xor (A(115) and B(90)) xor (A(116) and B(89)) xor (A(117) and B(88)) xor (A(118) and B(87)) xor (A(119) and B(86)) xor (A(120) and B(85)) xor (A(121) and B(84)) xor (A(122) and B(83)) xor (A(123) and B(82)) xor (A(124) and B(81)) xor (A(125) and B(80)) xor (A(126) and B(79)) xor (A(79) and B(127)) xor (A(80) and B(126)) xor (A(81) and B(125)) xor (A(82) and B(124)) xor (A(83) and B(123)) xor (A(84) and B(122)) xor (A(85) and B(121)) xor (A(86) and B(120)) xor (A(87) and B(119)) xor (A(88) and B(118)) xor (A(89) and B(117)) xor (A(90) and B(116)) xor (A(91) and B(115)) xor (A(92) and B(114)) xor (A(93) and B(113)) xor (A(94) and B(112)) xor (A(95) and B(111)) xor (A(96) and B(110)) xor (A(97) and B(109)) xor (A(98) and B(108)) xor (A(99) and B(107)) xor (A(100) and B(106)) xor (A(101) and B(105)) xor (A(102) and B(104)) xor (A(103) and B(103)) xor (A(104) and B(102)) xor (A(105) and B(101)) xor (A(106) and B(100)) xor (A(107) and B(99)) xor (A(108) and B(98)) xor (A(109) and B(97)) xor (A(110) and B(96)) xor (A(111) and B(95)) xor (A(112) and B(94)) xor (A(113) and B(93)) xor (A(114) and B(92)) xor (A(115) and B(91)) xor (A(116) and B(90)) xor (A(117) and B(89)) xor (A(118) and B(88)) xor (A(119) and B(87)) xor (A(120) and B(86)) xor (A(121) and B(85)) xor (A(122) and B(84)) xor (A(123) and B(83)) xor (A(124) and B(82)) xor (A(125) and B(81)) xor (A(126) and B(81));
    C(80)  <= (A(0) and B(80)) xor (A(1) and B(79)) xor (A(2) and B(78)) xor (A(3) and B(77)) xor (A(4) and B(76)) xor (A(5) and B(75)) xor (A(6) and B(74)) xor (A(7) and B(73)) xor (A(8) and B(72)) xor (A(9) and B(71)) xor (A(10) and B(70)) xor (A(11) and B(69)) xor (A(12) and B(68)) xor (A(13) and B(67)) xor (A(14) and B(66)) xor (A(15) and B(65)) xor (A(16) and B(64)) xor (A(17) and B(63)) xor (A(18) and B(62)) xor (A(19) and B(61)) xor (A(20) and B(60)) xor (A(21) and B(59)) xor (A(23) and B(58)) xor (A(23) and B(57)) xor (A(24) and B(56)) xor (A(25) and B(55)) xor (A(26) and B(54)) xor (A(27) and B(53)) xor (A(28) and B(52)) xor (A(29) and B(51)) xor (A(30) and B(50)) xor (A(31) and B(49)) xor (A(32) and B(48)) xor (A(33) and B(47)) xor (A(34) and B(46)) xor (A(35) and B(45)) xor (A(36) and B(44)) xor (A(37) and B(43)) xor (A(38) and B(42)) xor (A(39) and B(41)) xor (A(40) and B(40)) xor (A(41) and B(39)) xor (A(42) and B(38)) xor (A(43) and B(37)) xor (A(44) and B(36)) xor (A(45) and B(35)) xor (A(46) and B(34)) xor (A(47) and B(33)) xor (A(48) and B(32)) xor (A(49) and B(31)) xor (A(50) and B(30)) xor (A(51) and B(29)) xor (A(52) and B(28)) xor (A(53) and B(27)) xor (A(54) and B(26)) xor (A(55) and B(25)) xor (A(56) and B(24)) xor (A(57) and B(23)) xor (A(58) and B(23)) xor (A(59) and B(21)) xor (A(60) and B(20)) xor (A(61) and B(19)) xor (A(62) and B(18)) xor (A(63) and B(17)) xor (A(64) and B(16)) xor (A(65) and B(15)) xor (A(66) and B(14)) xor (A(67) and B(13)) xor (A(68) and B(12)) xor (A(69) and B(11)) xor (A(70) and B(10)) xor (A(71) and B(9)) xor (A(72) and B(8)) xor (A(73) and B(7)) xor (A(74) and B(6)) xor (A(75) and B(5)) xor (A(76) and B(4)) xor (A(77) and B(3)) xor (A(78) and B(2)) xor (A(79) and B(1)) xor (A(80) and B(0)) xor (A(73) and B(127)) xor (A(74) and B(126)) xor (A(75) and B(125)) xor (A(76) and B(124)) xor (A(77) and B(123)) xor (A(78) and B(122)) xor (A(79) and B(121)) xor (A(80) and B(120)) xor (A(81) and B(119)) xor (A(82) and B(118)) xor (A(83) and B(117)) xor (A(84) and B(116)) xor (A(85) and B(115)) xor (A(86) and B(114)) xor (A(87) and B(113)) xor (A(88) and B(112)) xor (A(89) and B(111)) xor (A(90) and B(110)) xor (A(91) and B(109)) xor (A(92) and B(108)) xor (A(93) and B(107)) xor (A(94) and B(106)) xor (A(95) and B(105)) xor (A(96) and B(104)) xor (A(97) and B(103)) xor (A(98) and B(102)) xor (A(99) and B(101)) xor (A(100) and B(100)) xor (A(101) and B(99)) xor (A(102) and B(98)) xor (A(103) and B(97)) xor (A(104) and B(96)) xor (A(105) and B(95)) xor (A(106) and B(94)) xor (A(107) and B(93)) xor (A(108) and B(92)) xor (A(109) and B(91)) xor (A(110) and B(90)) xor (A(111) and B(89)) xor (A(112) and B(88)) xor (A(113) and B(87)) xor (A(114) and B(86)) xor (A(115) and B(85)) xor (A(116) and B(84)) xor (A(117) and B(83)) xor (A(118) and B(82)) xor (A(119) and B(81)) xor (A(120) and B(80)) xor (A(121) and B(79)) xor (A(122) and B(78)) xor (A(123) and B(77)) xor (A(124) and B(76)) xor (A(125) and B(75)) xor (A(126) and B(74)) xor (A(78) and B(127)) xor (A(79) and B(126)) xor (A(80) and B(125)) xor (A(81) and B(124)) xor (A(82) and B(123)) xor (A(83) and B(122)) xor (A(84) and B(121)) xor (A(85) and B(120)) xor (A(86) and B(119)) xor (A(87) and B(118)) xor (A(88) and B(117)) xor (A(89) and B(116)) xor (A(90) and B(115)) xor (A(91) and B(114)) xor (A(92) and B(113)) xor (A(93) and B(112)) xor (A(94) and B(111)) xor (A(95) and B(110)) xor (A(96) and B(109)) xor (A(97) and B(108)) xor (A(98) and B(107)) xor (A(99) and B(106)) xor (A(100) and B(105)) xor (A(101) and B(104)) xor (A(102) and B(103)) xor (A(103) and B(102)) xor (A(104) and B(101)) xor (A(105) and B(100)) xor (A(106) and B(99)) xor (A(107) and B(98)) xor (A(108) and B(97)) xor (A(109) and B(96)) xor (A(110) and B(95)) xor (A(111) and B(94)) xor (A(112) and B(93)) xor (A(113) and B(92)) xor (A(114) and B(91)) xor (A(115) and B(90)) xor (A(116) and B(89)) xor (A(117) and B(88)) xor (A(118) and B(87)) xor (A(119) and B(86)) xor (A(120) and B(85)) xor (A(121) and B(84)) xor (A(122) and B(83)) xor (A(123) and B(82)) xor (A(124) and B(81)) xor (A(125) and B(80)) xor (A(126) and B(79)) xor (A(79) and B(127)) xor (A(80) and B(126)) xor (A(81) and B(125)) xor (A(82) and B(124)) xor (A(83) and B(123)) xor (A(84) and B(122)) xor (A(85) and B(121)) xor (A(86) and B(120)) xor (A(87) and B(119)) xor (A(88) and B(118)) xor (A(89) and B(117)) xor (A(90) and B(116)) xor (A(91) and B(115)) xor (A(92) and B(114)) xor (A(93) and B(113)) xor (A(94) and B(112)) xor (A(95) and B(111)) xor (A(96) and B(110)) xor (A(97) and B(109)) xor (A(98) and B(108)) xor (A(99) and B(107)) xor (A(100) and B(106)) xor (A(101) and B(105)) xor (A(102) and B(104)) xor (A(103) and B(103)) xor (A(104) and B(102)) xor (A(105) and B(101)) xor (A(106) and B(100)) xor (A(107) and B(99)) xor (A(108) and B(98)) xor (A(109) and B(97)) xor (A(110) and B(96)) xor (A(111) and B(95)) xor (A(112) and B(94)) xor (A(113) and B(93)) xor (A(114) and B(92)) xor (A(115) and B(91)) xor (A(116) and B(90)) xor (A(117) and B(89)) xor (A(118) and B(88)) xor (A(119) and B(87)) xor (A(120) and B(86)) xor (A(121) and B(85)) xor (A(122) and B(84)) xor (A(123) and B(83)) xor (A(124) and B(82)) xor (A(125) and B(81)) xor (A(126) and B(80)) xor (A(80) and B(127)) xor (A(81) and B(126)) xor (A(82) and B(125)) xor (A(83) and B(124)) xor (A(84) and B(123)) xor (A(85) and B(122)) xor (A(86) and B(121)) xor (A(87) and B(120)) xor (A(88) and B(119)) xor (A(89) and B(118)) xor (A(90) and B(117)) xor (A(91) and B(116)) xor (A(92) and B(115)) xor (A(93) and B(114)) xor (A(94) and B(113)) xor (A(95) and B(112)) xor (A(96) and B(111)) xor (A(97) and B(110)) xor (A(98) and B(109)) xor (A(99) and B(108)) xor (A(100) and B(107)) xor (A(101) and B(106)) xor (A(102) and B(105)) xor (A(103) and B(104)) xor (A(104) and B(103)) xor (A(105) and B(102)) xor (A(106) and B(101)) xor (A(107) and B(100)) xor (A(108) and B(99)) xor (A(109) and B(98)) xor (A(110) and B(97)) xor (A(111) and B(96)) xor (A(112) and B(95)) xor (A(113) and B(94)) xor (A(114) and B(93)) xor (A(115) and B(92)) xor (A(116) and B(91)) xor (A(117) and B(90)) xor (A(118) and B(89)) xor (A(119) and B(88)) xor (A(120) and B(87)) xor (A(121) and B(86)) xor (A(122) and B(85)) xor (A(123) and B(84)) xor (A(124) and B(83)) xor (A(125) and B(82)) xor (A(126) and B(82));
    C(81)  <= (A(0) and B(81)) xor (A(1) and B(80)) xor (A(2) and B(79)) xor (A(3) and B(78)) xor (A(4) and B(77)) xor (A(5) and B(76)) xor (A(6) and B(75)) xor (A(7) and B(74)) xor (A(8) and B(73)) xor (A(9) and B(72)) xor (A(10) and B(71)) xor (A(11) and B(70)) xor (A(12) and B(69)) xor (A(13) and B(68)) xor (A(14) and B(67)) xor (A(15) and B(66)) xor (A(16) and B(65)) xor (A(17) and B(64)) xor (A(18) and B(63)) xor (A(19) and B(62)) xor (A(20) and B(61)) xor (A(21) and B(60)) xor (A(23) and B(59)) xor (A(23) and B(58)) xor (A(24) and B(57)) xor (A(25) and B(56)) xor (A(26) and B(55)) xor (A(27) and B(54)) xor (A(28) and B(53)) xor (A(29) and B(52)) xor (A(30) and B(51)) xor (A(31) and B(50)) xor (A(32) and B(49)) xor (A(33) and B(48)) xor (A(34) and B(47)) xor (A(35) and B(46)) xor (A(36) and B(45)) xor (A(37) and B(44)) xor (A(38) and B(43)) xor (A(39) and B(42)) xor (A(40) and B(41)) xor (A(41) and B(40)) xor (A(42) and B(39)) xor (A(43) and B(38)) xor (A(44) and B(37)) xor (A(45) and B(36)) xor (A(46) and B(35)) xor (A(47) and B(34)) xor (A(48) and B(33)) xor (A(49) and B(32)) xor (A(50) and B(31)) xor (A(51) and B(30)) xor (A(52) and B(29)) xor (A(53) and B(28)) xor (A(54) and B(27)) xor (A(55) and B(26)) xor (A(56) and B(25)) xor (A(57) and B(24)) xor (A(58) and B(23)) xor (A(59) and B(23)) xor (A(60) and B(21)) xor (A(61) and B(20)) xor (A(62) and B(19)) xor (A(63) and B(18)) xor (A(64) and B(17)) xor (A(65) and B(16)) xor (A(66) and B(15)) xor (A(67) and B(14)) xor (A(68) and B(13)) xor (A(69) and B(12)) xor (A(70) and B(11)) xor (A(71) and B(10)) xor (A(72) and B(9)) xor (A(73) and B(8)) xor (A(74) and B(7)) xor (A(75) and B(6)) xor (A(76) and B(5)) xor (A(77) and B(4)) xor (A(78) and B(3)) xor (A(79) and B(2)) xor (A(80) and B(1)) xor (A(81) and B(0)) xor (A(74) and B(127)) xor (A(75) and B(126)) xor (A(76) and B(125)) xor (A(77) and B(124)) xor (A(78) and B(123)) xor (A(79) and B(122)) xor (A(80) and B(121)) xor (A(81) and B(120)) xor (A(82) and B(119)) xor (A(83) and B(118)) xor (A(84) and B(117)) xor (A(85) and B(116)) xor (A(86) and B(115)) xor (A(87) and B(114)) xor (A(88) and B(113)) xor (A(89) and B(112)) xor (A(90) and B(111)) xor (A(91) and B(110)) xor (A(92) and B(109)) xor (A(93) and B(108)) xor (A(94) and B(107)) xor (A(95) and B(106)) xor (A(96) and B(105)) xor (A(97) and B(104)) xor (A(98) and B(103)) xor (A(99) and B(102)) xor (A(100) and B(101)) xor (A(101) and B(100)) xor (A(102) and B(99)) xor (A(103) and B(98)) xor (A(104) and B(97)) xor (A(105) and B(96)) xor (A(106) and B(95)) xor (A(107) and B(94)) xor (A(108) and B(93)) xor (A(109) and B(92)) xor (A(110) and B(91)) xor (A(111) and B(90)) xor (A(112) and B(89)) xor (A(113) and B(88)) xor (A(114) and B(87)) xor (A(115) and B(86)) xor (A(116) and B(85)) xor (A(117) and B(84)) xor (A(118) and B(83)) xor (A(119) and B(82)) xor (A(120) and B(81)) xor (A(121) and B(80)) xor (A(122) and B(79)) xor (A(123) and B(78)) xor (A(124) and B(77)) xor (A(125) and B(76)) xor (A(126) and B(75)) xor (A(79) and B(127)) xor (A(80) and B(126)) xor (A(81) and B(125)) xor (A(82) and B(124)) xor (A(83) and B(123)) xor (A(84) and B(122)) xor (A(85) and B(121)) xor (A(86) and B(120)) xor (A(87) and B(119)) xor (A(88) and B(118)) xor (A(89) and B(117)) xor (A(90) and B(116)) xor (A(91) and B(115)) xor (A(92) and B(114)) xor (A(93) and B(113)) xor (A(94) and B(112)) xor (A(95) and B(111)) xor (A(96) and B(110)) xor (A(97) and B(109)) xor (A(98) and B(108)) xor (A(99) and B(107)) xor (A(100) and B(106)) xor (A(101) and B(105)) xor (A(102) and B(104)) xor (A(103) and B(103)) xor (A(104) and B(102)) xor (A(105) and B(101)) xor (A(106) and B(100)) xor (A(107) and B(99)) xor (A(108) and B(98)) xor (A(109) and B(97)) xor (A(110) and B(96)) xor (A(111) and B(95)) xor (A(112) and B(94)) xor (A(113) and B(93)) xor (A(114) and B(92)) xor (A(115) and B(91)) xor (A(116) and B(90)) xor (A(117) and B(89)) xor (A(118) and B(88)) xor (A(119) and B(87)) xor (A(120) and B(86)) xor (A(121) and B(85)) xor (A(122) and B(84)) xor (A(123) and B(83)) xor (A(124) and B(82)) xor (A(125) and B(81)) xor (A(126) and B(80)) xor (A(80) and B(127)) xor (A(81) and B(126)) xor (A(82) and B(125)) xor (A(83) and B(124)) xor (A(84) and B(123)) xor (A(85) and B(122)) xor (A(86) and B(121)) xor (A(87) and B(120)) xor (A(88) and B(119)) xor (A(89) and B(118)) xor (A(90) and B(117)) xor (A(91) and B(116)) xor (A(92) and B(115)) xor (A(93) and B(114)) xor (A(94) and B(113)) xor (A(95) and B(112)) xor (A(96) and B(111)) xor (A(97) and B(110)) xor (A(98) and B(109)) xor (A(99) and B(108)) xor (A(100) and B(107)) xor (A(101) and B(106)) xor (A(102) and B(105)) xor (A(103) and B(104)) xor (A(104) and B(103)) xor (A(105) and B(102)) xor (A(106) and B(101)) xor (A(107) and B(100)) xor (A(108) and B(99)) xor (A(109) and B(98)) xor (A(110) and B(97)) xor (A(111) and B(96)) xor (A(112) and B(95)) xor (A(113) and B(94)) xor (A(114) and B(93)) xor (A(115) and B(92)) xor (A(116) and B(91)) xor (A(117) and B(90)) xor (A(118) and B(89)) xor (A(119) and B(88)) xor (A(120) and B(87)) xor (A(121) and B(86)) xor (A(122) and B(85)) xor (A(123) and B(84)) xor (A(124) and B(83)) xor (A(125) and B(82)) xor (A(126) and B(81)) xor (A(81) and B(127)) xor (A(82) and B(126)) xor (A(83) and B(125)) xor (A(84) and B(124)) xor (A(85) and B(123)) xor (A(86) and B(122)) xor (A(87) and B(121)) xor (A(88) and B(120)) xor (A(89) and B(119)) xor (A(90) and B(118)) xor (A(91) and B(117)) xor (A(92) and B(116)) xor (A(93) and B(115)) xor (A(94) and B(114)) xor (A(95) and B(113)) xor (A(96) and B(112)) xor (A(97) and B(111)) xor (A(98) and B(110)) xor (A(99) and B(109)) xor (A(100) and B(108)) xor (A(101) and B(107)) xor (A(102) and B(106)) xor (A(103) and B(105)) xor (A(104) and B(104)) xor (A(105) and B(103)) xor (A(106) and B(102)) xor (A(107) and B(101)) xor (A(108) and B(100)) xor (A(109) and B(99)) xor (A(110) and B(98)) xor (A(111) and B(97)) xor (A(112) and B(96)) xor (A(113) and B(95)) xor (A(114) and B(94)) xor (A(115) and B(93)) xor (A(116) and B(92)) xor (A(117) and B(91)) xor (A(118) and B(90)) xor (A(119) and B(89)) xor (A(120) and B(88)) xor (A(121) and B(87)) xor (A(122) and B(86)) xor (A(123) and B(85)) xor (A(124) and B(84)) xor (A(125) and B(83)) xor (A(126) and B(83));
    C(82)  <= (A(0) and B(82)) xor (A(1) and B(81)) xor (A(2) and B(80)) xor (A(3) and B(79)) xor (A(4) and B(78)) xor (A(5) and B(77)) xor (A(6) and B(76)) xor (A(7) and B(75)) xor (A(8) and B(74)) xor (A(9) and B(73)) xor (A(10) and B(72)) xor (A(11) and B(71)) xor (A(12) and B(70)) xor (A(13) and B(69)) xor (A(14) and B(68)) xor (A(15) and B(67)) xor (A(16) and B(66)) xor (A(17) and B(65)) xor (A(18) and B(64)) xor (A(19) and B(63)) xor (A(20) and B(62)) xor (A(21) and B(61)) xor (A(23) and B(60)) xor (A(23) and B(59)) xor (A(24) and B(58)) xor (A(25) and B(57)) xor (A(26) and B(56)) xor (A(27) and B(55)) xor (A(28) and B(54)) xor (A(29) and B(53)) xor (A(30) and B(52)) xor (A(31) and B(51)) xor (A(32) and B(50)) xor (A(33) and B(49)) xor (A(34) and B(48)) xor (A(35) and B(47)) xor (A(36) and B(46)) xor (A(37) and B(45)) xor (A(38) and B(44)) xor (A(39) and B(43)) xor (A(40) and B(42)) xor (A(41) and B(41)) xor (A(42) and B(40)) xor (A(43) and B(39)) xor (A(44) and B(38)) xor (A(45) and B(37)) xor (A(46) and B(36)) xor (A(47) and B(35)) xor (A(48) and B(34)) xor (A(49) and B(33)) xor (A(50) and B(32)) xor (A(51) and B(31)) xor (A(52) and B(30)) xor (A(53) and B(29)) xor (A(54) and B(28)) xor (A(55) and B(27)) xor (A(56) and B(26)) xor (A(57) and B(25)) xor (A(58) and B(24)) xor (A(59) and B(23)) xor (A(60) and B(23)) xor (A(61) and B(21)) xor (A(62) and B(20)) xor (A(63) and B(19)) xor (A(64) and B(18)) xor (A(65) and B(17)) xor (A(66) and B(16)) xor (A(67) and B(15)) xor (A(68) and B(14)) xor (A(69) and B(13)) xor (A(70) and B(12)) xor (A(71) and B(11)) xor (A(72) and B(10)) xor (A(73) and B(9)) xor (A(74) and B(8)) xor (A(75) and B(7)) xor (A(76) and B(6)) xor (A(77) and B(5)) xor (A(78) and B(4)) xor (A(79) and B(3)) xor (A(80) and B(2)) xor (A(81) and B(1)) xor (A(82) and B(0)) xor (A(75) and B(127)) xor (A(76) and B(126)) xor (A(77) and B(125)) xor (A(78) and B(124)) xor (A(79) and B(123)) xor (A(80) and B(122)) xor (A(81) and B(121)) xor (A(82) and B(120)) xor (A(83) and B(119)) xor (A(84) and B(118)) xor (A(85) and B(117)) xor (A(86) and B(116)) xor (A(87) and B(115)) xor (A(88) and B(114)) xor (A(89) and B(113)) xor (A(90) and B(112)) xor (A(91) and B(111)) xor (A(92) and B(110)) xor (A(93) and B(109)) xor (A(94) and B(108)) xor (A(95) and B(107)) xor (A(96) and B(106)) xor (A(97) and B(105)) xor (A(98) and B(104)) xor (A(99) and B(103)) xor (A(100) and B(102)) xor (A(101) and B(101)) xor (A(102) and B(100)) xor (A(103) and B(99)) xor (A(104) and B(98)) xor (A(105) and B(97)) xor (A(106) and B(96)) xor (A(107) and B(95)) xor (A(108) and B(94)) xor (A(109) and B(93)) xor (A(110) and B(92)) xor (A(111) and B(91)) xor (A(112) and B(90)) xor (A(113) and B(89)) xor (A(114) and B(88)) xor (A(115) and B(87)) xor (A(116) and B(86)) xor (A(117) and B(85)) xor (A(118) and B(84)) xor (A(119) and B(83)) xor (A(120) and B(82)) xor (A(121) and B(81)) xor (A(122) and B(80)) xor (A(123) and B(79)) xor (A(124) and B(78)) xor (A(125) and B(77)) xor (A(126) and B(76)) xor (A(80) and B(127)) xor (A(81) and B(126)) xor (A(82) and B(125)) xor (A(83) and B(124)) xor (A(84) and B(123)) xor (A(85) and B(122)) xor (A(86) and B(121)) xor (A(87) and B(120)) xor (A(88) and B(119)) xor (A(89) and B(118)) xor (A(90) and B(117)) xor (A(91) and B(116)) xor (A(92) and B(115)) xor (A(93) and B(114)) xor (A(94) and B(113)) xor (A(95) and B(112)) xor (A(96) and B(111)) xor (A(97) and B(110)) xor (A(98) and B(109)) xor (A(99) and B(108)) xor (A(100) and B(107)) xor (A(101) and B(106)) xor (A(102) and B(105)) xor (A(103) and B(104)) xor (A(104) and B(103)) xor (A(105) and B(102)) xor (A(106) and B(101)) xor (A(107) and B(100)) xor (A(108) and B(99)) xor (A(109) and B(98)) xor (A(110) and B(97)) xor (A(111) and B(96)) xor (A(112) and B(95)) xor (A(113) and B(94)) xor (A(114) and B(93)) xor (A(115) and B(92)) xor (A(116) and B(91)) xor (A(117) and B(90)) xor (A(118) and B(89)) xor (A(119) and B(88)) xor (A(120) and B(87)) xor (A(121) and B(86)) xor (A(122) and B(85)) xor (A(123) and B(84)) xor (A(124) and B(83)) xor (A(125) and B(82)) xor (A(126) and B(81)) xor (A(81) and B(127)) xor (A(82) and B(126)) xor (A(83) and B(125)) xor (A(84) and B(124)) xor (A(85) and B(123)) xor (A(86) and B(122)) xor (A(87) and B(121)) xor (A(88) and B(120)) xor (A(89) and B(119)) xor (A(90) and B(118)) xor (A(91) and B(117)) xor (A(92) and B(116)) xor (A(93) and B(115)) xor (A(94) and B(114)) xor (A(95) and B(113)) xor (A(96) and B(112)) xor (A(97) and B(111)) xor (A(98) and B(110)) xor (A(99) and B(109)) xor (A(100) and B(108)) xor (A(101) and B(107)) xor (A(102) and B(106)) xor (A(103) and B(105)) xor (A(104) and B(104)) xor (A(105) and B(103)) xor (A(106) and B(102)) xor (A(107) and B(101)) xor (A(108) and B(100)) xor (A(109) and B(99)) xor (A(110) and B(98)) xor (A(111) and B(97)) xor (A(112) and B(96)) xor (A(113) and B(95)) xor (A(114) and B(94)) xor (A(115) and B(93)) xor (A(116) and B(92)) xor (A(117) and B(91)) xor (A(118) and B(90)) xor (A(119) and B(89)) xor (A(120) and B(88)) xor (A(121) and B(87)) xor (A(122) and B(86)) xor (A(123) and B(85)) xor (A(124) and B(84)) xor (A(125) and B(83)) xor (A(126) and B(82)) xor (A(82) and B(127)) xor (A(83) and B(126)) xor (A(84) and B(125)) xor (A(85) and B(124)) xor (A(86) and B(123)) xor (A(87) and B(122)) xor (A(88) and B(121)) xor (A(89) and B(120)) xor (A(90) and B(119)) xor (A(91) and B(118)) xor (A(92) and B(117)) xor (A(93) and B(116)) xor (A(94) and B(115)) xor (A(95) and B(114)) xor (A(96) and B(113)) xor (A(97) and B(112)) xor (A(98) and B(111)) xor (A(99) and B(110)) xor (A(100) and B(109)) xor (A(101) and B(108)) xor (A(102) and B(107)) xor (A(103) and B(106)) xor (A(104) and B(105)) xor (A(105) and B(104)) xor (A(106) and B(103)) xor (A(107) and B(102)) xor (A(108) and B(101)) xor (A(109) and B(100)) xor (A(110) and B(99)) xor (A(111) and B(98)) xor (A(112) and B(97)) xor (A(113) and B(96)) xor (A(114) and B(95)) xor (A(115) and B(94)) xor (A(116) and B(93)) xor (A(117) and B(92)) xor (A(118) and B(91)) xor (A(119) and B(90)) xor (A(120) and B(89)) xor (A(121) and B(88)) xor (A(122) and B(87)) xor (A(123) and B(86)) xor (A(124) and B(85)) xor (A(125) and B(84)) xor (A(126) and B(84));
    C(83)  <= (A(0) and B(83)) xor (A(1) and B(82)) xor (A(2) and B(81)) xor (A(3) and B(80)) xor (A(4) and B(79)) xor (A(5) and B(78)) xor (A(6) and B(77)) xor (A(7) and B(76)) xor (A(8) and B(75)) xor (A(9) and B(74)) xor (A(10) and B(73)) xor (A(11) and B(72)) xor (A(12) and B(71)) xor (A(13) and B(70)) xor (A(14) and B(69)) xor (A(15) and B(68)) xor (A(16) and B(67)) xor (A(17) and B(66)) xor (A(18) and B(65)) xor (A(19) and B(64)) xor (A(20) and B(63)) xor (A(21) and B(62)) xor (A(23) and B(61)) xor (A(23) and B(60)) xor (A(24) and B(59)) xor (A(25) and B(58)) xor (A(26) and B(57)) xor (A(27) and B(56)) xor (A(28) and B(55)) xor (A(29) and B(54)) xor (A(30) and B(53)) xor (A(31) and B(52)) xor (A(32) and B(51)) xor (A(33) and B(50)) xor (A(34) and B(49)) xor (A(35) and B(48)) xor (A(36) and B(47)) xor (A(37) and B(46)) xor (A(38) and B(45)) xor (A(39) and B(44)) xor (A(40) and B(43)) xor (A(41) and B(42)) xor (A(42) and B(41)) xor (A(43) and B(40)) xor (A(44) and B(39)) xor (A(45) and B(38)) xor (A(46) and B(37)) xor (A(47) and B(36)) xor (A(48) and B(35)) xor (A(49) and B(34)) xor (A(50) and B(33)) xor (A(51) and B(32)) xor (A(52) and B(31)) xor (A(53) and B(30)) xor (A(54) and B(29)) xor (A(55) and B(28)) xor (A(56) and B(27)) xor (A(57) and B(26)) xor (A(58) and B(25)) xor (A(59) and B(24)) xor (A(60) and B(23)) xor (A(61) and B(23)) xor (A(62) and B(21)) xor (A(63) and B(20)) xor (A(64) and B(19)) xor (A(65) and B(18)) xor (A(66) and B(17)) xor (A(67) and B(16)) xor (A(68) and B(15)) xor (A(69) and B(14)) xor (A(70) and B(13)) xor (A(71) and B(12)) xor (A(72) and B(11)) xor (A(73) and B(10)) xor (A(74) and B(9)) xor (A(75) and B(8)) xor (A(76) and B(7)) xor (A(77) and B(6)) xor (A(78) and B(5)) xor (A(79) and B(4)) xor (A(80) and B(3)) xor (A(81) and B(2)) xor (A(82) and B(1)) xor (A(83) and B(0)) xor (A(76) and B(127)) xor (A(77) and B(126)) xor (A(78) and B(125)) xor (A(79) and B(124)) xor (A(80) and B(123)) xor (A(81) and B(122)) xor (A(82) and B(121)) xor (A(83) and B(120)) xor (A(84) and B(119)) xor (A(85) and B(118)) xor (A(86) and B(117)) xor (A(87) and B(116)) xor (A(88) and B(115)) xor (A(89) and B(114)) xor (A(90) and B(113)) xor (A(91) and B(112)) xor (A(92) and B(111)) xor (A(93) and B(110)) xor (A(94) and B(109)) xor (A(95) and B(108)) xor (A(96) and B(107)) xor (A(97) and B(106)) xor (A(98) and B(105)) xor (A(99) and B(104)) xor (A(100) and B(103)) xor (A(101) and B(102)) xor (A(102) and B(101)) xor (A(103) and B(100)) xor (A(104) and B(99)) xor (A(105) and B(98)) xor (A(106) and B(97)) xor (A(107) and B(96)) xor (A(108) and B(95)) xor (A(109) and B(94)) xor (A(110) and B(93)) xor (A(111) and B(92)) xor (A(112) and B(91)) xor (A(113) and B(90)) xor (A(114) and B(89)) xor (A(115) and B(88)) xor (A(116) and B(87)) xor (A(117) and B(86)) xor (A(118) and B(85)) xor (A(119) and B(84)) xor (A(120) and B(83)) xor (A(121) and B(82)) xor (A(122) and B(81)) xor (A(123) and B(80)) xor (A(124) and B(79)) xor (A(125) and B(78)) xor (A(126) and B(77)) xor (A(81) and B(127)) xor (A(82) and B(126)) xor (A(83) and B(125)) xor (A(84) and B(124)) xor (A(85) and B(123)) xor (A(86) and B(122)) xor (A(87) and B(121)) xor (A(88) and B(120)) xor (A(89) and B(119)) xor (A(90) and B(118)) xor (A(91) and B(117)) xor (A(92) and B(116)) xor (A(93) and B(115)) xor (A(94) and B(114)) xor (A(95) and B(113)) xor (A(96) and B(112)) xor (A(97) and B(111)) xor (A(98) and B(110)) xor (A(99) and B(109)) xor (A(100) and B(108)) xor (A(101) and B(107)) xor (A(102) and B(106)) xor (A(103) and B(105)) xor (A(104) and B(104)) xor (A(105) and B(103)) xor (A(106) and B(102)) xor (A(107) and B(101)) xor (A(108) and B(100)) xor (A(109) and B(99)) xor (A(110) and B(98)) xor (A(111) and B(97)) xor (A(112) and B(96)) xor (A(113) and B(95)) xor (A(114) and B(94)) xor (A(115) and B(93)) xor (A(116) and B(92)) xor (A(117) and B(91)) xor (A(118) and B(90)) xor (A(119) and B(89)) xor (A(120) and B(88)) xor (A(121) and B(87)) xor (A(122) and B(86)) xor (A(123) and B(85)) xor (A(124) and B(84)) xor (A(125) and B(83)) xor (A(126) and B(82)) xor (A(82) and B(127)) xor (A(83) and B(126)) xor (A(84) and B(125)) xor (A(85) and B(124)) xor (A(86) and B(123)) xor (A(87) and B(122)) xor (A(88) and B(121)) xor (A(89) and B(120)) xor (A(90) and B(119)) xor (A(91) and B(118)) xor (A(92) and B(117)) xor (A(93) and B(116)) xor (A(94) and B(115)) xor (A(95) and B(114)) xor (A(96) and B(113)) xor (A(97) and B(112)) xor (A(98) and B(111)) xor (A(99) and B(110)) xor (A(100) and B(109)) xor (A(101) and B(108)) xor (A(102) and B(107)) xor (A(103) and B(106)) xor (A(104) and B(105)) xor (A(105) and B(104)) xor (A(106) and B(103)) xor (A(107) and B(102)) xor (A(108) and B(101)) xor (A(109) and B(100)) xor (A(110) and B(99)) xor (A(111) and B(98)) xor (A(112) and B(97)) xor (A(113) and B(96)) xor (A(114) and B(95)) xor (A(115) and B(94)) xor (A(116) and B(93)) xor (A(117) and B(92)) xor (A(118) and B(91)) xor (A(119) and B(90)) xor (A(120) and B(89)) xor (A(121) and B(88)) xor (A(122) and B(87)) xor (A(123) and B(86)) xor (A(124) and B(85)) xor (A(125) and B(84)) xor (A(126) and B(83)) xor (A(83) and B(127)) xor (A(84) and B(126)) xor (A(85) and B(125)) xor (A(86) and B(124)) xor (A(87) and B(123)) xor (A(88) and B(122)) xor (A(89) and B(121)) xor (A(90) and B(120)) xor (A(91) and B(119)) xor (A(92) and B(118)) xor (A(93) and B(117)) xor (A(94) and B(116)) xor (A(95) and B(115)) xor (A(96) and B(114)) xor (A(97) and B(113)) xor (A(98) and B(112)) xor (A(99) and B(111)) xor (A(100) and B(110)) xor (A(101) and B(109)) xor (A(102) and B(108)) xor (A(103) and B(107)) xor (A(104) and B(106)) xor (A(105) and B(105)) xor (A(106) and B(104)) xor (A(107) and B(103)) xor (A(108) and B(102)) xor (A(109) and B(101)) xor (A(110) and B(100)) xor (A(111) and B(99)) xor (A(112) and B(98)) xor (A(113) and B(97)) xor (A(114) and B(96)) xor (A(115) and B(95)) xor (A(116) and B(94)) xor (A(117) and B(93)) xor (A(118) and B(92)) xor (A(119) and B(91)) xor (A(120) and B(90)) xor (A(121) and B(89)) xor (A(122) and B(88)) xor (A(123) and B(87)) xor (A(124) and B(86)) xor (A(125) and B(85)) xor (A(126) and B(85));
    C(84)  <= (A(0) and B(84)) xor (A(1) and B(83)) xor (A(2) and B(82)) xor (A(3) and B(81)) xor (A(4) and B(80)) xor (A(5) and B(79)) xor (A(6) and B(78)) xor (A(7) and B(77)) xor (A(8) and B(76)) xor (A(9) and B(75)) xor (A(10) and B(74)) xor (A(11) and B(73)) xor (A(12) and B(72)) xor (A(13) and B(71)) xor (A(14) and B(70)) xor (A(15) and B(69)) xor (A(16) and B(68)) xor (A(17) and B(67)) xor (A(18) and B(66)) xor (A(19) and B(65)) xor (A(20) and B(64)) xor (A(21) and B(63)) xor (A(23) and B(62)) xor (A(23) and B(61)) xor (A(24) and B(60)) xor (A(25) and B(59)) xor (A(26) and B(58)) xor (A(27) and B(57)) xor (A(28) and B(56)) xor (A(29) and B(55)) xor (A(30) and B(54)) xor (A(31) and B(53)) xor (A(32) and B(52)) xor (A(33) and B(51)) xor (A(34) and B(50)) xor (A(35) and B(49)) xor (A(36) and B(48)) xor (A(37) and B(47)) xor (A(38) and B(46)) xor (A(39) and B(45)) xor (A(40) and B(44)) xor (A(41) and B(43)) xor (A(42) and B(42)) xor (A(43) and B(41)) xor (A(44) and B(40)) xor (A(45) and B(39)) xor (A(46) and B(38)) xor (A(47) and B(37)) xor (A(48) and B(36)) xor (A(49) and B(35)) xor (A(50) and B(34)) xor (A(51) and B(33)) xor (A(52) and B(32)) xor (A(53) and B(31)) xor (A(54) and B(30)) xor (A(55) and B(29)) xor (A(56) and B(28)) xor (A(57) and B(27)) xor (A(58) and B(26)) xor (A(59) and B(25)) xor (A(60) and B(24)) xor (A(61) and B(23)) xor (A(62) and B(23)) xor (A(63) and B(21)) xor (A(64) and B(20)) xor (A(65) and B(19)) xor (A(66) and B(18)) xor (A(67) and B(17)) xor (A(68) and B(16)) xor (A(69) and B(15)) xor (A(70) and B(14)) xor (A(71) and B(13)) xor (A(72) and B(12)) xor (A(73) and B(11)) xor (A(74) and B(10)) xor (A(75) and B(9)) xor (A(76) and B(8)) xor (A(77) and B(7)) xor (A(78) and B(6)) xor (A(79) and B(5)) xor (A(80) and B(4)) xor (A(81) and B(3)) xor (A(82) and B(2)) xor (A(83) and B(1)) xor (A(84) and B(0)) xor (A(77) and B(127)) xor (A(78) and B(126)) xor (A(79) and B(125)) xor (A(80) and B(124)) xor (A(81) and B(123)) xor (A(82) and B(122)) xor (A(83) and B(121)) xor (A(84) and B(120)) xor (A(85) and B(119)) xor (A(86) and B(118)) xor (A(87) and B(117)) xor (A(88) and B(116)) xor (A(89) and B(115)) xor (A(90) and B(114)) xor (A(91) and B(113)) xor (A(92) and B(112)) xor (A(93) and B(111)) xor (A(94) and B(110)) xor (A(95) and B(109)) xor (A(96) and B(108)) xor (A(97) and B(107)) xor (A(98) and B(106)) xor (A(99) and B(105)) xor (A(100) and B(104)) xor (A(101) and B(103)) xor (A(102) and B(102)) xor (A(103) and B(101)) xor (A(104) and B(100)) xor (A(105) and B(99)) xor (A(106) and B(98)) xor (A(107) and B(97)) xor (A(108) and B(96)) xor (A(109) and B(95)) xor (A(110) and B(94)) xor (A(111) and B(93)) xor (A(112) and B(92)) xor (A(113) and B(91)) xor (A(114) and B(90)) xor (A(115) and B(89)) xor (A(116) and B(88)) xor (A(117) and B(87)) xor (A(118) and B(86)) xor (A(119) and B(85)) xor (A(120) and B(84)) xor (A(121) and B(83)) xor (A(122) and B(82)) xor (A(123) and B(81)) xor (A(124) and B(80)) xor (A(125) and B(79)) xor (A(126) and B(78)) xor (A(82) and B(127)) xor (A(83) and B(126)) xor (A(84) and B(125)) xor (A(85) and B(124)) xor (A(86) and B(123)) xor (A(87) and B(122)) xor (A(88) and B(121)) xor (A(89) and B(120)) xor (A(90) and B(119)) xor (A(91) and B(118)) xor (A(92) and B(117)) xor (A(93) and B(116)) xor (A(94) and B(115)) xor (A(95) and B(114)) xor (A(96) and B(113)) xor (A(97) and B(112)) xor (A(98) and B(111)) xor (A(99) and B(110)) xor (A(100) and B(109)) xor (A(101) and B(108)) xor (A(102) and B(107)) xor (A(103) and B(106)) xor (A(104) and B(105)) xor (A(105) and B(104)) xor (A(106) and B(103)) xor (A(107) and B(102)) xor (A(108) and B(101)) xor (A(109) and B(100)) xor (A(110) and B(99)) xor (A(111) and B(98)) xor (A(112) and B(97)) xor (A(113) and B(96)) xor (A(114) and B(95)) xor (A(115) and B(94)) xor (A(116) and B(93)) xor (A(117) and B(92)) xor (A(118) and B(91)) xor (A(119) and B(90)) xor (A(120) and B(89)) xor (A(121) and B(88)) xor (A(122) and B(87)) xor (A(123) and B(86)) xor (A(124) and B(85)) xor (A(125) and B(84)) xor (A(126) and B(83)) xor (A(83) and B(127)) xor (A(84) and B(126)) xor (A(85) and B(125)) xor (A(86) and B(124)) xor (A(87) and B(123)) xor (A(88) and B(122)) xor (A(89) and B(121)) xor (A(90) and B(120)) xor (A(91) and B(119)) xor (A(92) and B(118)) xor (A(93) and B(117)) xor (A(94) and B(116)) xor (A(95) and B(115)) xor (A(96) and B(114)) xor (A(97) and B(113)) xor (A(98) and B(112)) xor (A(99) and B(111)) xor (A(100) and B(110)) xor (A(101) and B(109)) xor (A(102) and B(108)) xor (A(103) and B(107)) xor (A(104) and B(106)) xor (A(105) and B(105)) xor (A(106) and B(104)) xor (A(107) and B(103)) xor (A(108) and B(102)) xor (A(109) and B(101)) xor (A(110) and B(100)) xor (A(111) and B(99)) xor (A(112) and B(98)) xor (A(113) and B(97)) xor (A(114) and B(96)) xor (A(115) and B(95)) xor (A(116) and B(94)) xor (A(117) and B(93)) xor (A(118) and B(92)) xor (A(119) and B(91)) xor (A(120) and B(90)) xor (A(121) and B(89)) xor (A(122) and B(88)) xor (A(123) and B(87)) xor (A(124) and B(86)) xor (A(125) and B(85)) xor (A(126) and B(84)) xor (A(84) and B(127)) xor (A(85) and B(126)) xor (A(86) and B(125)) xor (A(87) and B(124)) xor (A(88) and B(123)) xor (A(89) and B(122)) xor (A(90) and B(121)) xor (A(91) and B(120)) xor (A(92) and B(119)) xor (A(93) and B(118)) xor (A(94) and B(117)) xor (A(95) and B(116)) xor (A(96) and B(115)) xor (A(97) and B(114)) xor (A(98) and B(113)) xor (A(99) and B(112)) xor (A(100) and B(111)) xor (A(101) and B(110)) xor (A(102) and B(109)) xor (A(103) and B(108)) xor (A(104) and B(107)) xor (A(105) and B(106)) xor (A(106) and B(105)) xor (A(107) and B(104)) xor (A(108) and B(103)) xor (A(109) and B(102)) xor (A(110) and B(101)) xor (A(111) and B(100)) xor (A(112) and B(99)) xor (A(113) and B(98)) xor (A(114) and B(97)) xor (A(115) and B(96)) xor (A(116) and B(95)) xor (A(117) and B(94)) xor (A(118) and B(93)) xor (A(119) and B(92)) xor (A(120) and B(91)) xor (A(121) and B(90)) xor (A(122) and B(89)) xor (A(123) and B(88)) xor (A(124) and B(87)) xor (A(125) and B(86)) xor (A(126) and B(86));
    C(85)  <= (A(0) and B(85)) xor (A(1) and B(84)) xor (A(2) and B(83)) xor (A(3) and B(82)) xor (A(4) and B(81)) xor (A(5) and B(80)) xor (A(6) and B(79)) xor (A(7) and B(78)) xor (A(8) and B(77)) xor (A(9) and B(76)) xor (A(10) and B(75)) xor (A(11) and B(74)) xor (A(12) and B(73)) xor (A(13) and B(72)) xor (A(14) and B(71)) xor (A(15) and B(70)) xor (A(16) and B(69)) xor (A(17) and B(68)) xor (A(18) and B(67)) xor (A(19) and B(66)) xor (A(20) and B(65)) xor (A(21) and B(64)) xor (A(23) and B(63)) xor (A(23) and B(62)) xor (A(24) and B(61)) xor (A(25) and B(60)) xor (A(26) and B(59)) xor (A(27) and B(58)) xor (A(28) and B(57)) xor (A(29) and B(56)) xor (A(30) and B(55)) xor (A(31) and B(54)) xor (A(32) and B(53)) xor (A(33) and B(52)) xor (A(34) and B(51)) xor (A(35) and B(50)) xor (A(36) and B(49)) xor (A(37) and B(48)) xor (A(38) and B(47)) xor (A(39) and B(46)) xor (A(40) and B(45)) xor (A(41) and B(44)) xor (A(42) and B(43)) xor (A(43) and B(42)) xor (A(44) and B(41)) xor (A(45) and B(40)) xor (A(46) and B(39)) xor (A(47) and B(38)) xor (A(48) and B(37)) xor (A(49) and B(36)) xor (A(50) and B(35)) xor (A(51) and B(34)) xor (A(52) and B(33)) xor (A(53) and B(32)) xor (A(54) and B(31)) xor (A(55) and B(30)) xor (A(56) and B(29)) xor (A(57) and B(28)) xor (A(58) and B(27)) xor (A(59) and B(26)) xor (A(60) and B(25)) xor (A(61) and B(24)) xor (A(62) and B(23)) xor (A(63) and B(23)) xor (A(64) and B(21)) xor (A(65) and B(20)) xor (A(66) and B(19)) xor (A(67) and B(18)) xor (A(68) and B(17)) xor (A(69) and B(16)) xor (A(70) and B(15)) xor (A(71) and B(14)) xor (A(72) and B(13)) xor (A(73) and B(12)) xor (A(74) and B(11)) xor (A(75) and B(10)) xor (A(76) and B(9)) xor (A(77) and B(8)) xor (A(78) and B(7)) xor (A(79) and B(6)) xor (A(80) and B(5)) xor (A(81) and B(4)) xor (A(82) and B(3)) xor (A(83) and B(2)) xor (A(84) and B(1)) xor (A(85) and B(0)) xor (A(78) and B(127)) xor (A(79) and B(126)) xor (A(80) and B(125)) xor (A(81) and B(124)) xor (A(82) and B(123)) xor (A(83) and B(122)) xor (A(84) and B(121)) xor (A(85) and B(120)) xor (A(86) and B(119)) xor (A(87) and B(118)) xor (A(88) and B(117)) xor (A(89) and B(116)) xor (A(90) and B(115)) xor (A(91) and B(114)) xor (A(92) and B(113)) xor (A(93) and B(112)) xor (A(94) and B(111)) xor (A(95) and B(110)) xor (A(96) and B(109)) xor (A(97) and B(108)) xor (A(98) and B(107)) xor (A(99) and B(106)) xor (A(100) and B(105)) xor (A(101) and B(104)) xor (A(102) and B(103)) xor (A(103) and B(102)) xor (A(104) and B(101)) xor (A(105) and B(100)) xor (A(106) and B(99)) xor (A(107) and B(98)) xor (A(108) and B(97)) xor (A(109) and B(96)) xor (A(110) and B(95)) xor (A(111) and B(94)) xor (A(112) and B(93)) xor (A(113) and B(92)) xor (A(114) and B(91)) xor (A(115) and B(90)) xor (A(116) and B(89)) xor (A(117) and B(88)) xor (A(118) and B(87)) xor (A(119) and B(86)) xor (A(120) and B(85)) xor (A(121) and B(84)) xor (A(122) and B(83)) xor (A(123) and B(82)) xor (A(124) and B(81)) xor (A(125) and B(80)) xor (A(126) and B(79)) xor (A(83) and B(127)) xor (A(84) and B(126)) xor (A(85) and B(125)) xor (A(86) and B(124)) xor (A(87) and B(123)) xor (A(88) and B(122)) xor (A(89) and B(121)) xor (A(90) and B(120)) xor (A(91) and B(119)) xor (A(92) and B(118)) xor (A(93) and B(117)) xor (A(94) and B(116)) xor (A(95) and B(115)) xor (A(96) and B(114)) xor (A(97) and B(113)) xor (A(98) and B(112)) xor (A(99) and B(111)) xor (A(100) and B(110)) xor (A(101) and B(109)) xor (A(102) and B(108)) xor (A(103) and B(107)) xor (A(104) and B(106)) xor (A(105) and B(105)) xor (A(106) and B(104)) xor (A(107) and B(103)) xor (A(108) and B(102)) xor (A(109) and B(101)) xor (A(110) and B(100)) xor (A(111) and B(99)) xor (A(112) and B(98)) xor (A(113) and B(97)) xor (A(114) and B(96)) xor (A(115) and B(95)) xor (A(116) and B(94)) xor (A(117) and B(93)) xor (A(118) and B(92)) xor (A(119) and B(91)) xor (A(120) and B(90)) xor (A(121) and B(89)) xor (A(122) and B(88)) xor (A(123) and B(87)) xor (A(124) and B(86)) xor (A(125) and B(85)) xor (A(126) and B(84)) xor (A(84) and B(127)) xor (A(85) and B(126)) xor (A(86) and B(125)) xor (A(87) and B(124)) xor (A(88) and B(123)) xor (A(89) and B(122)) xor (A(90) and B(121)) xor (A(91) and B(120)) xor (A(92) and B(119)) xor (A(93) and B(118)) xor (A(94) and B(117)) xor (A(95) and B(116)) xor (A(96) and B(115)) xor (A(97) and B(114)) xor (A(98) and B(113)) xor (A(99) and B(112)) xor (A(100) and B(111)) xor (A(101) and B(110)) xor (A(102) and B(109)) xor (A(103) and B(108)) xor (A(104) and B(107)) xor (A(105) and B(106)) xor (A(106) and B(105)) xor (A(107) and B(104)) xor (A(108) and B(103)) xor (A(109) and B(102)) xor (A(110) and B(101)) xor (A(111) and B(100)) xor (A(112) and B(99)) xor (A(113) and B(98)) xor (A(114) and B(97)) xor (A(115) and B(96)) xor (A(116) and B(95)) xor (A(117) and B(94)) xor (A(118) and B(93)) xor (A(119) and B(92)) xor (A(120) and B(91)) xor (A(121) and B(90)) xor (A(122) and B(89)) xor (A(123) and B(88)) xor (A(124) and B(87)) xor (A(125) and B(86)) xor (A(126) and B(85)) xor (A(85) and B(127)) xor (A(86) and B(126)) xor (A(87) and B(125)) xor (A(88) and B(124)) xor (A(89) and B(123)) xor (A(90) and B(122)) xor (A(91) and B(121)) xor (A(92) and B(120)) xor (A(93) and B(119)) xor (A(94) and B(118)) xor (A(95) and B(117)) xor (A(96) and B(116)) xor (A(97) and B(115)) xor (A(98) and B(114)) xor (A(99) and B(113)) xor (A(100) and B(112)) xor (A(101) and B(111)) xor (A(102) and B(110)) xor (A(103) and B(109)) xor (A(104) and B(108)) xor (A(105) and B(107)) xor (A(106) and B(106)) xor (A(107) and B(105)) xor (A(108) and B(104)) xor (A(109) and B(103)) xor (A(110) and B(102)) xor (A(111) and B(101)) xor (A(112) and B(100)) xor (A(113) and B(99)) xor (A(114) and B(98)) xor (A(115) and B(97)) xor (A(116) and B(96)) xor (A(117) and B(95)) xor (A(118) and B(94)) xor (A(119) and B(93)) xor (A(120) and B(92)) xor (A(121) and B(91)) xor (A(122) and B(90)) xor (A(123) and B(89)) xor (A(124) and B(88)) xor (A(125) and B(87)) xor (A(126) and B(87));
    C(86)  <= (A(0) and B(86)) xor (A(1) and B(85)) xor (A(2) and B(84)) xor (A(3) and B(83)) xor (A(4) and B(82)) xor (A(5) and B(81)) xor (A(6) and B(80)) xor (A(7) and B(79)) xor (A(8) and B(78)) xor (A(9) and B(77)) xor (A(10) and B(76)) xor (A(11) and B(75)) xor (A(12) and B(74)) xor (A(13) and B(73)) xor (A(14) and B(72)) xor (A(15) and B(71)) xor (A(16) and B(70)) xor (A(17) and B(69)) xor (A(18) and B(68)) xor (A(19) and B(67)) xor (A(20) and B(66)) xor (A(21) and B(65)) xor (A(23) and B(64)) xor (A(23) and B(63)) xor (A(24) and B(62)) xor (A(25) and B(61)) xor (A(26) and B(60)) xor (A(27) and B(59)) xor (A(28) and B(58)) xor (A(29) and B(57)) xor (A(30) and B(56)) xor (A(31) and B(55)) xor (A(32) and B(54)) xor (A(33) and B(53)) xor (A(34) and B(52)) xor (A(35) and B(51)) xor (A(36) and B(50)) xor (A(37) and B(49)) xor (A(38) and B(48)) xor (A(39) and B(47)) xor (A(40) and B(46)) xor (A(41) and B(45)) xor (A(42) and B(44)) xor (A(43) and B(43)) xor (A(44) and B(42)) xor (A(45) and B(41)) xor (A(46) and B(40)) xor (A(47) and B(39)) xor (A(48) and B(38)) xor (A(49) and B(37)) xor (A(50) and B(36)) xor (A(51) and B(35)) xor (A(52) and B(34)) xor (A(53) and B(33)) xor (A(54) and B(32)) xor (A(55) and B(31)) xor (A(56) and B(30)) xor (A(57) and B(29)) xor (A(58) and B(28)) xor (A(59) and B(27)) xor (A(60) and B(26)) xor (A(61) and B(25)) xor (A(62) and B(24)) xor (A(63) and B(23)) xor (A(64) and B(23)) xor (A(65) and B(21)) xor (A(66) and B(20)) xor (A(67) and B(19)) xor (A(68) and B(18)) xor (A(69) and B(17)) xor (A(70) and B(16)) xor (A(71) and B(15)) xor (A(72) and B(14)) xor (A(73) and B(13)) xor (A(74) and B(12)) xor (A(75) and B(11)) xor (A(76) and B(10)) xor (A(77) and B(9)) xor (A(78) and B(8)) xor (A(79) and B(7)) xor (A(80) and B(6)) xor (A(81) and B(5)) xor (A(82) and B(4)) xor (A(83) and B(3)) xor (A(84) and B(2)) xor (A(85) and B(1)) xor (A(86) and B(0)) xor (A(79) and B(127)) xor (A(80) and B(126)) xor (A(81) and B(125)) xor (A(82) and B(124)) xor (A(83) and B(123)) xor (A(84) and B(122)) xor (A(85) and B(121)) xor (A(86) and B(120)) xor (A(87) and B(119)) xor (A(88) and B(118)) xor (A(89) and B(117)) xor (A(90) and B(116)) xor (A(91) and B(115)) xor (A(92) and B(114)) xor (A(93) and B(113)) xor (A(94) and B(112)) xor (A(95) and B(111)) xor (A(96) and B(110)) xor (A(97) and B(109)) xor (A(98) and B(108)) xor (A(99) and B(107)) xor (A(100) and B(106)) xor (A(101) and B(105)) xor (A(102) and B(104)) xor (A(103) and B(103)) xor (A(104) and B(102)) xor (A(105) and B(101)) xor (A(106) and B(100)) xor (A(107) and B(99)) xor (A(108) and B(98)) xor (A(109) and B(97)) xor (A(110) and B(96)) xor (A(111) and B(95)) xor (A(112) and B(94)) xor (A(113) and B(93)) xor (A(114) and B(92)) xor (A(115) and B(91)) xor (A(116) and B(90)) xor (A(117) and B(89)) xor (A(118) and B(88)) xor (A(119) and B(87)) xor (A(120) and B(86)) xor (A(121) and B(85)) xor (A(122) and B(84)) xor (A(123) and B(83)) xor (A(124) and B(82)) xor (A(125) and B(81)) xor (A(126) and B(80)) xor (A(84) and B(127)) xor (A(85) and B(126)) xor (A(86) and B(125)) xor (A(87) and B(124)) xor (A(88) and B(123)) xor (A(89) and B(122)) xor (A(90) and B(121)) xor (A(91) and B(120)) xor (A(92) and B(119)) xor (A(93) and B(118)) xor (A(94) and B(117)) xor (A(95) and B(116)) xor (A(96) and B(115)) xor (A(97) and B(114)) xor (A(98) and B(113)) xor (A(99) and B(112)) xor (A(100) and B(111)) xor (A(101) and B(110)) xor (A(102) and B(109)) xor (A(103) and B(108)) xor (A(104) and B(107)) xor (A(105) and B(106)) xor (A(106) and B(105)) xor (A(107) and B(104)) xor (A(108) and B(103)) xor (A(109) and B(102)) xor (A(110) and B(101)) xor (A(111) and B(100)) xor (A(112) and B(99)) xor (A(113) and B(98)) xor (A(114) and B(97)) xor (A(115) and B(96)) xor (A(116) and B(95)) xor (A(117) and B(94)) xor (A(118) and B(93)) xor (A(119) and B(92)) xor (A(120) and B(91)) xor (A(121) and B(90)) xor (A(122) and B(89)) xor (A(123) and B(88)) xor (A(124) and B(87)) xor (A(125) and B(86)) xor (A(126) and B(85)) xor (A(85) and B(127)) xor (A(86) and B(126)) xor (A(87) and B(125)) xor (A(88) and B(124)) xor (A(89) and B(123)) xor (A(90) and B(122)) xor (A(91) and B(121)) xor (A(92) and B(120)) xor (A(93) and B(119)) xor (A(94) and B(118)) xor (A(95) and B(117)) xor (A(96) and B(116)) xor (A(97) and B(115)) xor (A(98) and B(114)) xor (A(99) and B(113)) xor (A(100) and B(112)) xor (A(101) and B(111)) xor (A(102) and B(110)) xor (A(103) and B(109)) xor (A(104) and B(108)) xor (A(105) and B(107)) xor (A(106) and B(106)) xor (A(107) and B(105)) xor (A(108) and B(104)) xor (A(109) and B(103)) xor (A(110) and B(102)) xor (A(111) and B(101)) xor (A(112) and B(100)) xor (A(113) and B(99)) xor (A(114) and B(98)) xor (A(115) and B(97)) xor (A(116) and B(96)) xor (A(117) and B(95)) xor (A(118) and B(94)) xor (A(119) and B(93)) xor (A(120) and B(92)) xor (A(121) and B(91)) xor (A(122) and B(90)) xor (A(123) and B(89)) xor (A(124) and B(88)) xor (A(125) and B(87)) xor (A(126) and B(86)) xor (A(86) and B(127)) xor (A(87) and B(126)) xor (A(88) and B(125)) xor (A(89) and B(124)) xor (A(90) and B(123)) xor (A(91) and B(122)) xor (A(92) and B(121)) xor (A(93) and B(120)) xor (A(94) and B(119)) xor (A(95) and B(118)) xor (A(96) and B(117)) xor (A(97) and B(116)) xor (A(98) and B(115)) xor (A(99) and B(114)) xor (A(100) and B(113)) xor (A(101) and B(112)) xor (A(102) and B(111)) xor (A(103) and B(110)) xor (A(104) and B(109)) xor (A(105) and B(108)) xor (A(106) and B(107)) xor (A(107) and B(106)) xor (A(108) and B(105)) xor (A(109) and B(104)) xor (A(110) and B(103)) xor (A(111) and B(102)) xor (A(112) and B(101)) xor (A(113) and B(100)) xor (A(114) and B(99)) xor (A(115) and B(98)) xor (A(116) and B(97)) xor (A(117) and B(96)) xor (A(118) and B(95)) xor (A(119) and B(94)) xor (A(120) and B(93)) xor (A(121) and B(92)) xor (A(122) and B(91)) xor (A(123) and B(90)) xor (A(124) and B(89)) xor (A(125) and B(88)) xor (A(126) and B(88));
    C(87)  <= (A(0) and B(87)) xor (A(1) and B(86)) xor (A(2) and B(85)) xor (A(3) and B(84)) xor (A(4) and B(83)) xor (A(5) and B(82)) xor (A(6) and B(81)) xor (A(7) and B(80)) xor (A(8) and B(79)) xor (A(9) and B(78)) xor (A(10) and B(77)) xor (A(11) and B(76)) xor (A(12) and B(75)) xor (A(13) and B(74)) xor (A(14) and B(73)) xor (A(15) and B(72)) xor (A(16) and B(71)) xor (A(17) and B(70)) xor (A(18) and B(69)) xor (A(19) and B(68)) xor (A(20) and B(67)) xor (A(21) and B(66)) xor (A(23) and B(65)) xor (A(23) and B(64)) xor (A(24) and B(63)) xor (A(25) and B(62)) xor (A(26) and B(61)) xor (A(27) and B(60)) xor (A(28) and B(59)) xor (A(29) and B(58)) xor (A(30) and B(57)) xor (A(31) and B(56)) xor (A(32) and B(55)) xor (A(33) and B(54)) xor (A(34) and B(53)) xor (A(35) and B(52)) xor (A(36) and B(51)) xor (A(37) and B(50)) xor (A(38) and B(49)) xor (A(39) and B(48)) xor (A(40) and B(47)) xor (A(41) and B(46)) xor (A(42) and B(45)) xor (A(43) and B(44)) xor (A(44) and B(43)) xor (A(45) and B(42)) xor (A(46) and B(41)) xor (A(47) and B(40)) xor (A(48) and B(39)) xor (A(49) and B(38)) xor (A(50) and B(37)) xor (A(51) and B(36)) xor (A(52) and B(35)) xor (A(53) and B(34)) xor (A(54) and B(33)) xor (A(55) and B(32)) xor (A(56) and B(31)) xor (A(57) and B(30)) xor (A(58) and B(29)) xor (A(59) and B(28)) xor (A(60) and B(27)) xor (A(61) and B(26)) xor (A(62) and B(25)) xor (A(63) and B(24)) xor (A(64) and B(23)) xor (A(65) and B(23)) xor (A(66) and B(21)) xor (A(67) and B(20)) xor (A(68) and B(19)) xor (A(69) and B(18)) xor (A(70) and B(17)) xor (A(71) and B(16)) xor (A(72) and B(15)) xor (A(73) and B(14)) xor (A(74) and B(13)) xor (A(75) and B(12)) xor (A(76) and B(11)) xor (A(77) and B(10)) xor (A(78) and B(9)) xor (A(79) and B(8)) xor (A(80) and B(7)) xor (A(81) and B(6)) xor (A(82) and B(5)) xor (A(83) and B(4)) xor (A(84) and B(3)) xor (A(85) and B(2)) xor (A(86) and B(1)) xor (A(87) and B(0)) xor (A(80) and B(127)) xor (A(81) and B(126)) xor (A(82) and B(125)) xor (A(83) and B(124)) xor (A(84) and B(123)) xor (A(85) and B(122)) xor (A(86) and B(121)) xor (A(87) and B(120)) xor (A(88) and B(119)) xor (A(89) and B(118)) xor (A(90) and B(117)) xor (A(91) and B(116)) xor (A(92) and B(115)) xor (A(93) and B(114)) xor (A(94) and B(113)) xor (A(95) and B(112)) xor (A(96) and B(111)) xor (A(97) and B(110)) xor (A(98) and B(109)) xor (A(99) and B(108)) xor (A(100) and B(107)) xor (A(101) and B(106)) xor (A(102) and B(105)) xor (A(103) and B(104)) xor (A(104) and B(103)) xor (A(105) and B(102)) xor (A(106) and B(101)) xor (A(107) and B(100)) xor (A(108) and B(99)) xor (A(109) and B(98)) xor (A(110) and B(97)) xor (A(111) and B(96)) xor (A(112) and B(95)) xor (A(113) and B(94)) xor (A(114) and B(93)) xor (A(115) and B(92)) xor (A(116) and B(91)) xor (A(117) and B(90)) xor (A(118) and B(89)) xor (A(119) and B(88)) xor (A(120) and B(87)) xor (A(121) and B(86)) xor (A(122) and B(85)) xor (A(123) and B(84)) xor (A(124) and B(83)) xor (A(125) and B(82)) xor (A(126) and B(81)) xor (A(85) and B(127)) xor (A(86) and B(126)) xor (A(87) and B(125)) xor (A(88) and B(124)) xor (A(89) and B(123)) xor (A(90) and B(122)) xor (A(91) and B(121)) xor (A(92) and B(120)) xor (A(93) and B(119)) xor (A(94) and B(118)) xor (A(95) and B(117)) xor (A(96) and B(116)) xor (A(97) and B(115)) xor (A(98) and B(114)) xor (A(99) and B(113)) xor (A(100) and B(112)) xor (A(101) and B(111)) xor (A(102) and B(110)) xor (A(103) and B(109)) xor (A(104) and B(108)) xor (A(105) and B(107)) xor (A(106) and B(106)) xor (A(107) and B(105)) xor (A(108) and B(104)) xor (A(109) and B(103)) xor (A(110) and B(102)) xor (A(111) and B(101)) xor (A(112) and B(100)) xor (A(113) and B(99)) xor (A(114) and B(98)) xor (A(115) and B(97)) xor (A(116) and B(96)) xor (A(117) and B(95)) xor (A(118) and B(94)) xor (A(119) and B(93)) xor (A(120) and B(92)) xor (A(121) and B(91)) xor (A(122) and B(90)) xor (A(123) and B(89)) xor (A(124) and B(88)) xor (A(125) and B(87)) xor (A(126) and B(86)) xor (A(86) and B(127)) xor (A(87) and B(126)) xor (A(88) and B(125)) xor (A(89) and B(124)) xor (A(90) and B(123)) xor (A(91) and B(122)) xor (A(92) and B(121)) xor (A(93) and B(120)) xor (A(94) and B(119)) xor (A(95) and B(118)) xor (A(96) and B(117)) xor (A(97) and B(116)) xor (A(98) and B(115)) xor (A(99) and B(114)) xor (A(100) and B(113)) xor (A(101) and B(112)) xor (A(102) and B(111)) xor (A(103) and B(110)) xor (A(104) and B(109)) xor (A(105) and B(108)) xor (A(106) and B(107)) xor (A(107) and B(106)) xor (A(108) and B(105)) xor (A(109) and B(104)) xor (A(110) and B(103)) xor (A(111) and B(102)) xor (A(112) and B(101)) xor (A(113) and B(100)) xor (A(114) and B(99)) xor (A(115) and B(98)) xor (A(116) and B(97)) xor (A(117) and B(96)) xor (A(118) and B(95)) xor (A(119) and B(94)) xor (A(120) and B(93)) xor (A(121) and B(92)) xor (A(122) and B(91)) xor (A(123) and B(90)) xor (A(124) and B(89)) xor (A(125) and B(88)) xor (A(126) and B(87)) xor (A(87) and B(127)) xor (A(88) and B(126)) xor (A(89) and B(125)) xor (A(90) and B(124)) xor (A(91) and B(123)) xor (A(92) and B(122)) xor (A(93) and B(121)) xor (A(94) and B(120)) xor (A(95) and B(119)) xor (A(96) and B(118)) xor (A(97) and B(117)) xor (A(98) and B(116)) xor (A(99) and B(115)) xor (A(100) and B(114)) xor (A(101) and B(113)) xor (A(102) and B(112)) xor (A(103) and B(111)) xor (A(104) and B(110)) xor (A(105) and B(109)) xor (A(106) and B(108)) xor (A(107) and B(107)) xor (A(108) and B(106)) xor (A(109) and B(105)) xor (A(110) and B(104)) xor (A(111) and B(103)) xor (A(112) and B(102)) xor (A(113) and B(101)) xor (A(114) and B(100)) xor (A(115) and B(99)) xor (A(116) and B(98)) xor (A(117) and B(97)) xor (A(118) and B(96)) xor (A(119) and B(95)) xor (A(120) and B(94)) xor (A(121) and B(93)) xor (A(122) and B(92)) xor (A(123) and B(91)) xor (A(124) and B(90)) xor (A(125) and B(89)) xor (A(126) and B(89));
    C(88)  <= (A(0) and B(88)) xor (A(1) and B(87)) xor (A(2) and B(86)) xor (A(3) and B(85)) xor (A(4) and B(84)) xor (A(5) and B(83)) xor (A(6) and B(82)) xor (A(7) and B(81)) xor (A(8) and B(80)) xor (A(9) and B(79)) xor (A(10) and B(78)) xor (A(11) and B(77)) xor (A(12) and B(76)) xor (A(13) and B(75)) xor (A(14) and B(74)) xor (A(15) and B(73)) xor (A(16) and B(72)) xor (A(17) and B(71)) xor (A(18) and B(70)) xor (A(19) and B(69)) xor (A(20) and B(68)) xor (A(21) and B(67)) xor (A(23) and B(66)) xor (A(23) and B(65)) xor (A(24) and B(64)) xor (A(25) and B(63)) xor (A(26) and B(62)) xor (A(27) and B(61)) xor (A(28) and B(60)) xor (A(29) and B(59)) xor (A(30) and B(58)) xor (A(31) and B(57)) xor (A(32) and B(56)) xor (A(33) and B(55)) xor (A(34) and B(54)) xor (A(35) and B(53)) xor (A(36) and B(52)) xor (A(37) and B(51)) xor (A(38) and B(50)) xor (A(39) and B(49)) xor (A(40) and B(48)) xor (A(41) and B(47)) xor (A(42) and B(46)) xor (A(43) and B(45)) xor (A(44) and B(44)) xor (A(45) and B(43)) xor (A(46) and B(42)) xor (A(47) and B(41)) xor (A(48) and B(40)) xor (A(49) and B(39)) xor (A(50) and B(38)) xor (A(51) and B(37)) xor (A(52) and B(36)) xor (A(53) and B(35)) xor (A(54) and B(34)) xor (A(55) and B(33)) xor (A(56) and B(32)) xor (A(57) and B(31)) xor (A(58) and B(30)) xor (A(59) and B(29)) xor (A(60) and B(28)) xor (A(61) and B(27)) xor (A(62) and B(26)) xor (A(63) and B(25)) xor (A(64) and B(24)) xor (A(65) and B(23)) xor (A(66) and B(23)) xor (A(67) and B(21)) xor (A(68) and B(20)) xor (A(69) and B(19)) xor (A(70) and B(18)) xor (A(71) and B(17)) xor (A(72) and B(16)) xor (A(73) and B(15)) xor (A(74) and B(14)) xor (A(75) and B(13)) xor (A(76) and B(12)) xor (A(77) and B(11)) xor (A(78) and B(10)) xor (A(79) and B(9)) xor (A(80) and B(8)) xor (A(81) and B(7)) xor (A(82) and B(6)) xor (A(83) and B(5)) xor (A(84) and B(4)) xor (A(85) and B(3)) xor (A(86) and B(2)) xor (A(87) and B(1)) xor (A(88) and B(0)) xor (A(81) and B(127)) xor (A(82) and B(126)) xor (A(83) and B(125)) xor (A(84) and B(124)) xor (A(85) and B(123)) xor (A(86) and B(122)) xor (A(87) and B(121)) xor (A(88) and B(120)) xor (A(89) and B(119)) xor (A(90) and B(118)) xor (A(91) and B(117)) xor (A(92) and B(116)) xor (A(93) and B(115)) xor (A(94) and B(114)) xor (A(95) and B(113)) xor (A(96) and B(112)) xor (A(97) and B(111)) xor (A(98) and B(110)) xor (A(99) and B(109)) xor (A(100) and B(108)) xor (A(101) and B(107)) xor (A(102) and B(106)) xor (A(103) and B(105)) xor (A(104) and B(104)) xor (A(105) and B(103)) xor (A(106) and B(102)) xor (A(107) and B(101)) xor (A(108) and B(100)) xor (A(109) and B(99)) xor (A(110) and B(98)) xor (A(111) and B(97)) xor (A(112) and B(96)) xor (A(113) and B(95)) xor (A(114) and B(94)) xor (A(115) and B(93)) xor (A(116) and B(92)) xor (A(117) and B(91)) xor (A(118) and B(90)) xor (A(119) and B(89)) xor (A(120) and B(88)) xor (A(121) and B(87)) xor (A(122) and B(86)) xor (A(123) and B(85)) xor (A(124) and B(84)) xor (A(125) and B(83)) xor (A(126) and B(82)) xor (A(86) and B(127)) xor (A(87) and B(126)) xor (A(88) and B(125)) xor (A(89) and B(124)) xor (A(90) and B(123)) xor (A(91) and B(122)) xor (A(92) and B(121)) xor (A(93) and B(120)) xor (A(94) and B(119)) xor (A(95) and B(118)) xor (A(96) and B(117)) xor (A(97) and B(116)) xor (A(98) and B(115)) xor (A(99) and B(114)) xor (A(100) and B(113)) xor (A(101) and B(112)) xor (A(102) and B(111)) xor (A(103) and B(110)) xor (A(104) and B(109)) xor (A(105) and B(108)) xor (A(106) and B(107)) xor (A(107) and B(106)) xor (A(108) and B(105)) xor (A(109) and B(104)) xor (A(110) and B(103)) xor (A(111) and B(102)) xor (A(112) and B(101)) xor (A(113) and B(100)) xor (A(114) and B(99)) xor (A(115) and B(98)) xor (A(116) and B(97)) xor (A(117) and B(96)) xor (A(118) and B(95)) xor (A(119) and B(94)) xor (A(120) and B(93)) xor (A(121) and B(92)) xor (A(122) and B(91)) xor (A(123) and B(90)) xor (A(124) and B(89)) xor (A(125) and B(88)) xor (A(126) and B(87)) xor (A(87) and B(127)) xor (A(88) and B(126)) xor (A(89) and B(125)) xor (A(90) and B(124)) xor (A(91) and B(123)) xor (A(92) and B(122)) xor (A(93) and B(121)) xor (A(94) and B(120)) xor (A(95) and B(119)) xor (A(96) and B(118)) xor (A(97) and B(117)) xor (A(98) and B(116)) xor (A(99) and B(115)) xor (A(100) and B(114)) xor (A(101) and B(113)) xor (A(102) and B(112)) xor (A(103) and B(111)) xor (A(104) and B(110)) xor (A(105) and B(109)) xor (A(106) and B(108)) xor (A(107) and B(107)) xor (A(108) and B(106)) xor (A(109) and B(105)) xor (A(110) and B(104)) xor (A(111) and B(103)) xor (A(112) and B(102)) xor (A(113) and B(101)) xor (A(114) and B(100)) xor (A(115) and B(99)) xor (A(116) and B(98)) xor (A(117) and B(97)) xor (A(118) and B(96)) xor (A(119) and B(95)) xor (A(120) and B(94)) xor (A(121) and B(93)) xor (A(122) and B(92)) xor (A(123) and B(91)) xor (A(124) and B(90)) xor (A(125) and B(89)) xor (A(126) and B(88)) xor (A(88) and B(127)) xor (A(89) and B(126)) xor (A(90) and B(125)) xor (A(91) and B(124)) xor (A(92) and B(123)) xor (A(93) and B(122)) xor (A(94) and B(121)) xor (A(95) and B(120)) xor (A(96) and B(119)) xor (A(97) and B(118)) xor (A(98) and B(117)) xor (A(99) and B(116)) xor (A(100) and B(115)) xor (A(101) and B(114)) xor (A(102) and B(113)) xor (A(103) and B(112)) xor (A(104) and B(111)) xor (A(105) and B(110)) xor (A(106) and B(109)) xor (A(107) and B(108)) xor (A(108) and B(107)) xor (A(109) and B(106)) xor (A(110) and B(105)) xor (A(111) and B(104)) xor (A(112) and B(103)) xor (A(113) and B(102)) xor (A(114) and B(101)) xor (A(115) and B(100)) xor (A(116) and B(99)) xor (A(117) and B(98)) xor (A(118) and B(97)) xor (A(119) and B(96)) xor (A(120) and B(95)) xor (A(121) and B(94)) xor (A(122) and B(93)) xor (A(123) and B(92)) xor (A(124) and B(91)) xor (A(125) and B(90)) xor (A(126) and B(90));
    C(89)  <= (A(0) and B(89)) xor (A(1) and B(88)) xor (A(2) and B(87)) xor (A(3) and B(86)) xor (A(4) and B(85)) xor (A(5) and B(84)) xor (A(6) and B(83)) xor (A(7) and B(82)) xor (A(8) and B(81)) xor (A(9) and B(80)) xor (A(10) and B(79)) xor (A(11) and B(78)) xor (A(12) and B(77)) xor (A(13) and B(76)) xor (A(14) and B(75)) xor (A(15) and B(74)) xor (A(16) and B(73)) xor (A(17) and B(72)) xor (A(18) and B(71)) xor (A(19) and B(70)) xor (A(20) and B(69)) xor (A(21) and B(68)) xor (A(23) and B(67)) xor (A(23) and B(66)) xor (A(24) and B(65)) xor (A(25) and B(64)) xor (A(26) and B(63)) xor (A(27) and B(62)) xor (A(28) and B(61)) xor (A(29) and B(60)) xor (A(30) and B(59)) xor (A(31) and B(58)) xor (A(32) and B(57)) xor (A(33) and B(56)) xor (A(34) and B(55)) xor (A(35) and B(54)) xor (A(36) and B(53)) xor (A(37) and B(52)) xor (A(38) and B(51)) xor (A(39) and B(50)) xor (A(40) and B(49)) xor (A(41) and B(48)) xor (A(42) and B(47)) xor (A(43) and B(46)) xor (A(44) and B(45)) xor (A(45) and B(44)) xor (A(46) and B(43)) xor (A(47) and B(42)) xor (A(48) and B(41)) xor (A(49) and B(40)) xor (A(50) and B(39)) xor (A(51) and B(38)) xor (A(52) and B(37)) xor (A(53) and B(36)) xor (A(54) and B(35)) xor (A(55) and B(34)) xor (A(56) and B(33)) xor (A(57) and B(32)) xor (A(58) and B(31)) xor (A(59) and B(30)) xor (A(60) and B(29)) xor (A(61) and B(28)) xor (A(62) and B(27)) xor (A(63) and B(26)) xor (A(64) and B(25)) xor (A(65) and B(24)) xor (A(66) and B(23)) xor (A(67) and B(23)) xor (A(68) and B(21)) xor (A(69) and B(20)) xor (A(70) and B(19)) xor (A(71) and B(18)) xor (A(72) and B(17)) xor (A(73) and B(16)) xor (A(74) and B(15)) xor (A(75) and B(14)) xor (A(76) and B(13)) xor (A(77) and B(12)) xor (A(78) and B(11)) xor (A(79) and B(10)) xor (A(80) and B(9)) xor (A(81) and B(8)) xor (A(82) and B(7)) xor (A(83) and B(6)) xor (A(84) and B(5)) xor (A(85) and B(4)) xor (A(86) and B(3)) xor (A(87) and B(2)) xor (A(88) and B(1)) xor (A(89) and B(0)) xor (A(82) and B(127)) xor (A(83) and B(126)) xor (A(84) and B(125)) xor (A(85) and B(124)) xor (A(86) and B(123)) xor (A(87) and B(122)) xor (A(88) and B(121)) xor (A(89) and B(120)) xor (A(90) and B(119)) xor (A(91) and B(118)) xor (A(92) and B(117)) xor (A(93) and B(116)) xor (A(94) and B(115)) xor (A(95) and B(114)) xor (A(96) and B(113)) xor (A(97) and B(112)) xor (A(98) and B(111)) xor (A(99) and B(110)) xor (A(100) and B(109)) xor (A(101) and B(108)) xor (A(102) and B(107)) xor (A(103) and B(106)) xor (A(104) and B(105)) xor (A(105) and B(104)) xor (A(106) and B(103)) xor (A(107) and B(102)) xor (A(108) and B(101)) xor (A(109) and B(100)) xor (A(110) and B(99)) xor (A(111) and B(98)) xor (A(112) and B(97)) xor (A(113) and B(96)) xor (A(114) and B(95)) xor (A(115) and B(94)) xor (A(116) and B(93)) xor (A(117) and B(92)) xor (A(118) and B(91)) xor (A(119) and B(90)) xor (A(120) and B(89)) xor (A(121) and B(88)) xor (A(122) and B(87)) xor (A(123) and B(86)) xor (A(124) and B(85)) xor (A(125) and B(84)) xor (A(126) and B(83)) xor (A(87) and B(127)) xor (A(88) and B(126)) xor (A(89) and B(125)) xor (A(90) and B(124)) xor (A(91) and B(123)) xor (A(92) and B(122)) xor (A(93) and B(121)) xor (A(94) and B(120)) xor (A(95) and B(119)) xor (A(96) and B(118)) xor (A(97) and B(117)) xor (A(98) and B(116)) xor (A(99) and B(115)) xor (A(100) and B(114)) xor (A(101) and B(113)) xor (A(102) and B(112)) xor (A(103) and B(111)) xor (A(104) and B(110)) xor (A(105) and B(109)) xor (A(106) and B(108)) xor (A(107) and B(107)) xor (A(108) and B(106)) xor (A(109) and B(105)) xor (A(110) and B(104)) xor (A(111) and B(103)) xor (A(112) and B(102)) xor (A(113) and B(101)) xor (A(114) and B(100)) xor (A(115) and B(99)) xor (A(116) and B(98)) xor (A(117) and B(97)) xor (A(118) and B(96)) xor (A(119) and B(95)) xor (A(120) and B(94)) xor (A(121) and B(93)) xor (A(122) and B(92)) xor (A(123) and B(91)) xor (A(124) and B(90)) xor (A(125) and B(89)) xor (A(126) and B(88)) xor (A(88) and B(127)) xor (A(89) and B(126)) xor (A(90) and B(125)) xor (A(91) and B(124)) xor (A(92) and B(123)) xor (A(93) and B(122)) xor (A(94) and B(121)) xor (A(95) and B(120)) xor (A(96) and B(119)) xor (A(97) and B(118)) xor (A(98) and B(117)) xor (A(99) and B(116)) xor (A(100) and B(115)) xor (A(101) and B(114)) xor (A(102) and B(113)) xor (A(103) and B(112)) xor (A(104) and B(111)) xor (A(105) and B(110)) xor (A(106) and B(109)) xor (A(107) and B(108)) xor (A(108) and B(107)) xor (A(109) and B(106)) xor (A(110) and B(105)) xor (A(111) and B(104)) xor (A(112) and B(103)) xor (A(113) and B(102)) xor (A(114) and B(101)) xor (A(115) and B(100)) xor (A(116) and B(99)) xor (A(117) and B(98)) xor (A(118) and B(97)) xor (A(119) and B(96)) xor (A(120) and B(95)) xor (A(121) and B(94)) xor (A(122) and B(93)) xor (A(123) and B(92)) xor (A(124) and B(91)) xor (A(125) and B(90)) xor (A(126) and B(89)) xor (A(89) and B(127)) xor (A(90) and B(126)) xor (A(91) and B(125)) xor (A(92) and B(124)) xor (A(93) and B(123)) xor (A(94) and B(122)) xor (A(95) and B(121)) xor (A(96) and B(120)) xor (A(97) and B(119)) xor (A(98) and B(118)) xor (A(99) and B(117)) xor (A(100) and B(116)) xor (A(101) and B(115)) xor (A(102) and B(114)) xor (A(103) and B(113)) xor (A(104) and B(112)) xor (A(105) and B(111)) xor (A(106) and B(110)) xor (A(107) and B(109)) xor (A(108) and B(108)) xor (A(109) and B(107)) xor (A(110) and B(106)) xor (A(111) and B(105)) xor (A(112) and B(104)) xor (A(113) and B(103)) xor (A(114) and B(102)) xor (A(115) and B(101)) xor (A(116) and B(100)) xor (A(117) and B(99)) xor (A(118) and B(98)) xor (A(119) and B(97)) xor (A(120) and B(96)) xor (A(121) and B(95)) xor (A(122) and B(94)) xor (A(123) and B(93)) xor (A(124) and B(92)) xor (A(125) and B(91)) xor (A(126) and B(91));
    C(90)  <= (A(0) and B(90)) xor (A(1) and B(89)) xor (A(2) and B(88)) xor (A(3) and B(87)) xor (A(4) and B(86)) xor (A(5) and B(85)) xor (A(6) and B(84)) xor (A(7) and B(83)) xor (A(8) and B(82)) xor (A(9) and B(81)) xor (A(10) and B(80)) xor (A(11) and B(79)) xor (A(12) and B(78)) xor (A(13) and B(77)) xor (A(14) and B(76)) xor (A(15) and B(75)) xor (A(16) and B(74)) xor (A(17) and B(73)) xor (A(18) and B(72)) xor (A(19) and B(71)) xor (A(20) and B(70)) xor (A(21) and B(69)) xor (A(23) and B(68)) xor (A(23) and B(67)) xor (A(24) and B(66)) xor (A(25) and B(65)) xor (A(26) and B(64)) xor (A(27) and B(63)) xor (A(28) and B(62)) xor (A(29) and B(61)) xor (A(30) and B(60)) xor (A(31) and B(59)) xor (A(32) and B(58)) xor (A(33) and B(57)) xor (A(34) and B(56)) xor (A(35) and B(55)) xor (A(36) and B(54)) xor (A(37) and B(53)) xor (A(38) and B(52)) xor (A(39) and B(51)) xor (A(40) and B(50)) xor (A(41) and B(49)) xor (A(42) and B(48)) xor (A(43) and B(47)) xor (A(44) and B(46)) xor (A(45) and B(45)) xor (A(46) and B(44)) xor (A(47) and B(43)) xor (A(48) and B(42)) xor (A(49) and B(41)) xor (A(50) and B(40)) xor (A(51) and B(39)) xor (A(52) and B(38)) xor (A(53) and B(37)) xor (A(54) and B(36)) xor (A(55) and B(35)) xor (A(56) and B(34)) xor (A(57) and B(33)) xor (A(58) and B(32)) xor (A(59) and B(31)) xor (A(60) and B(30)) xor (A(61) and B(29)) xor (A(62) and B(28)) xor (A(63) and B(27)) xor (A(64) and B(26)) xor (A(65) and B(25)) xor (A(66) and B(24)) xor (A(67) and B(23)) xor (A(68) and B(23)) xor (A(69) and B(21)) xor (A(70) and B(20)) xor (A(71) and B(19)) xor (A(72) and B(18)) xor (A(73) and B(17)) xor (A(74) and B(16)) xor (A(75) and B(15)) xor (A(76) and B(14)) xor (A(77) and B(13)) xor (A(78) and B(12)) xor (A(79) and B(11)) xor (A(80) and B(10)) xor (A(81) and B(9)) xor (A(82) and B(8)) xor (A(83) and B(7)) xor (A(84) and B(6)) xor (A(85) and B(5)) xor (A(86) and B(4)) xor (A(87) and B(3)) xor (A(88) and B(2)) xor (A(89) and B(1)) xor (A(90) and B(0)) xor (A(83) and B(127)) xor (A(84) and B(126)) xor (A(85) and B(125)) xor (A(86) and B(124)) xor (A(87) and B(123)) xor (A(88) and B(122)) xor (A(89) and B(121)) xor (A(90) and B(120)) xor (A(91) and B(119)) xor (A(92) and B(118)) xor (A(93) and B(117)) xor (A(94) and B(116)) xor (A(95) and B(115)) xor (A(96) and B(114)) xor (A(97) and B(113)) xor (A(98) and B(112)) xor (A(99) and B(111)) xor (A(100) and B(110)) xor (A(101) and B(109)) xor (A(102) and B(108)) xor (A(103) and B(107)) xor (A(104) and B(106)) xor (A(105) and B(105)) xor (A(106) and B(104)) xor (A(107) and B(103)) xor (A(108) and B(102)) xor (A(109) and B(101)) xor (A(110) and B(100)) xor (A(111) and B(99)) xor (A(112) and B(98)) xor (A(113) and B(97)) xor (A(114) and B(96)) xor (A(115) and B(95)) xor (A(116) and B(94)) xor (A(117) and B(93)) xor (A(118) and B(92)) xor (A(119) and B(91)) xor (A(120) and B(90)) xor (A(121) and B(89)) xor (A(122) and B(88)) xor (A(123) and B(87)) xor (A(124) and B(86)) xor (A(125) and B(85)) xor (A(126) and B(84)) xor (A(88) and B(127)) xor (A(89) and B(126)) xor (A(90) and B(125)) xor (A(91) and B(124)) xor (A(92) and B(123)) xor (A(93) and B(122)) xor (A(94) and B(121)) xor (A(95) and B(120)) xor (A(96) and B(119)) xor (A(97) and B(118)) xor (A(98) and B(117)) xor (A(99) and B(116)) xor (A(100) and B(115)) xor (A(101) and B(114)) xor (A(102) and B(113)) xor (A(103) and B(112)) xor (A(104) and B(111)) xor (A(105) and B(110)) xor (A(106) and B(109)) xor (A(107) and B(108)) xor (A(108) and B(107)) xor (A(109) and B(106)) xor (A(110) and B(105)) xor (A(111) and B(104)) xor (A(112) and B(103)) xor (A(113) and B(102)) xor (A(114) and B(101)) xor (A(115) and B(100)) xor (A(116) and B(99)) xor (A(117) and B(98)) xor (A(118) and B(97)) xor (A(119) and B(96)) xor (A(120) and B(95)) xor (A(121) and B(94)) xor (A(122) and B(93)) xor (A(123) and B(92)) xor (A(124) and B(91)) xor (A(125) and B(90)) xor (A(126) and B(89)) xor (A(89) and B(127)) xor (A(90) and B(126)) xor (A(91) and B(125)) xor (A(92) and B(124)) xor (A(93) and B(123)) xor (A(94) and B(122)) xor (A(95) and B(121)) xor (A(96) and B(120)) xor (A(97) and B(119)) xor (A(98) and B(118)) xor (A(99) and B(117)) xor (A(100) and B(116)) xor (A(101) and B(115)) xor (A(102) and B(114)) xor (A(103) and B(113)) xor (A(104) and B(112)) xor (A(105) and B(111)) xor (A(106) and B(110)) xor (A(107) and B(109)) xor (A(108) and B(108)) xor (A(109) and B(107)) xor (A(110) and B(106)) xor (A(111) and B(105)) xor (A(112) and B(104)) xor (A(113) and B(103)) xor (A(114) and B(102)) xor (A(115) and B(101)) xor (A(116) and B(100)) xor (A(117) and B(99)) xor (A(118) and B(98)) xor (A(119) and B(97)) xor (A(120) and B(96)) xor (A(121) and B(95)) xor (A(122) and B(94)) xor (A(123) and B(93)) xor (A(124) and B(92)) xor (A(125) and B(91)) xor (A(126) and B(90)) xor (A(90) and B(127)) xor (A(91) and B(126)) xor (A(92) and B(125)) xor (A(93) and B(124)) xor (A(94) and B(123)) xor (A(95) and B(122)) xor (A(96) and B(121)) xor (A(97) and B(120)) xor (A(98) and B(119)) xor (A(99) and B(118)) xor (A(100) and B(117)) xor (A(101) and B(116)) xor (A(102) and B(115)) xor (A(103) and B(114)) xor (A(104) and B(113)) xor (A(105) and B(112)) xor (A(106) and B(111)) xor (A(107) and B(110)) xor (A(108) and B(109)) xor (A(109) and B(108)) xor (A(110) and B(107)) xor (A(111) and B(106)) xor (A(112) and B(105)) xor (A(113) and B(104)) xor (A(114) and B(103)) xor (A(115) and B(102)) xor (A(116) and B(101)) xor (A(117) and B(100)) xor (A(118) and B(99)) xor (A(119) and B(98)) xor (A(120) and B(97)) xor (A(121) and B(96)) xor (A(122) and B(95)) xor (A(123) and B(94)) xor (A(124) and B(93)) xor (A(125) and B(92)) xor (A(126) and B(92));
    C(91)  <= (A(0) and B(91)) xor (A(1) and B(90)) xor (A(2) and B(89)) xor (A(3) and B(88)) xor (A(4) and B(87)) xor (A(5) and B(86)) xor (A(6) and B(85)) xor (A(7) and B(84)) xor (A(8) and B(83)) xor (A(9) and B(82)) xor (A(10) and B(81)) xor (A(11) and B(80)) xor (A(12) and B(79)) xor (A(13) and B(78)) xor (A(14) and B(77)) xor (A(15) and B(76)) xor (A(16) and B(75)) xor (A(17) and B(74)) xor (A(18) and B(73)) xor (A(19) and B(72)) xor (A(20) and B(71)) xor (A(21) and B(70)) xor (A(23) and B(69)) xor (A(23) and B(68)) xor (A(24) and B(67)) xor (A(25) and B(66)) xor (A(26) and B(65)) xor (A(27) and B(64)) xor (A(28) and B(63)) xor (A(29) and B(62)) xor (A(30) and B(61)) xor (A(31) and B(60)) xor (A(32) and B(59)) xor (A(33) and B(58)) xor (A(34) and B(57)) xor (A(35) and B(56)) xor (A(36) and B(55)) xor (A(37) and B(54)) xor (A(38) and B(53)) xor (A(39) and B(52)) xor (A(40) and B(51)) xor (A(41) and B(50)) xor (A(42) and B(49)) xor (A(43) and B(48)) xor (A(44) and B(47)) xor (A(45) and B(46)) xor (A(46) and B(45)) xor (A(47) and B(44)) xor (A(48) and B(43)) xor (A(49) and B(42)) xor (A(50) and B(41)) xor (A(51) and B(40)) xor (A(52) and B(39)) xor (A(53) and B(38)) xor (A(54) and B(37)) xor (A(55) and B(36)) xor (A(56) and B(35)) xor (A(57) and B(34)) xor (A(58) and B(33)) xor (A(59) and B(32)) xor (A(60) and B(31)) xor (A(61) and B(30)) xor (A(62) and B(29)) xor (A(63) and B(28)) xor (A(64) and B(27)) xor (A(65) and B(26)) xor (A(66) and B(25)) xor (A(67) and B(24)) xor (A(68) and B(23)) xor (A(69) and B(23)) xor (A(70) and B(21)) xor (A(71) and B(20)) xor (A(72) and B(19)) xor (A(73) and B(18)) xor (A(74) and B(17)) xor (A(75) and B(16)) xor (A(76) and B(15)) xor (A(77) and B(14)) xor (A(78) and B(13)) xor (A(79) and B(12)) xor (A(80) and B(11)) xor (A(81) and B(10)) xor (A(82) and B(9)) xor (A(83) and B(8)) xor (A(84) and B(7)) xor (A(85) and B(6)) xor (A(86) and B(5)) xor (A(87) and B(4)) xor (A(88) and B(3)) xor (A(89) and B(2)) xor (A(90) and B(1)) xor (A(91) and B(0)) xor (A(84) and B(127)) xor (A(85) and B(126)) xor (A(86) and B(125)) xor (A(87) and B(124)) xor (A(88) and B(123)) xor (A(89) and B(122)) xor (A(90) and B(121)) xor (A(91) and B(120)) xor (A(92) and B(119)) xor (A(93) and B(118)) xor (A(94) and B(117)) xor (A(95) and B(116)) xor (A(96) and B(115)) xor (A(97) and B(114)) xor (A(98) and B(113)) xor (A(99) and B(112)) xor (A(100) and B(111)) xor (A(101) and B(110)) xor (A(102) and B(109)) xor (A(103) and B(108)) xor (A(104) and B(107)) xor (A(105) and B(106)) xor (A(106) and B(105)) xor (A(107) and B(104)) xor (A(108) and B(103)) xor (A(109) and B(102)) xor (A(110) and B(101)) xor (A(111) and B(100)) xor (A(112) and B(99)) xor (A(113) and B(98)) xor (A(114) and B(97)) xor (A(115) and B(96)) xor (A(116) and B(95)) xor (A(117) and B(94)) xor (A(118) and B(93)) xor (A(119) and B(92)) xor (A(120) and B(91)) xor (A(121) and B(90)) xor (A(122) and B(89)) xor (A(123) and B(88)) xor (A(124) and B(87)) xor (A(125) and B(86)) xor (A(126) and B(85)) xor (A(89) and B(127)) xor (A(90) and B(126)) xor (A(91) and B(125)) xor (A(92) and B(124)) xor (A(93) and B(123)) xor (A(94) and B(122)) xor (A(95) and B(121)) xor (A(96) and B(120)) xor (A(97) and B(119)) xor (A(98) and B(118)) xor (A(99) and B(117)) xor (A(100) and B(116)) xor (A(101) and B(115)) xor (A(102) and B(114)) xor (A(103) and B(113)) xor (A(104) and B(112)) xor (A(105) and B(111)) xor (A(106) and B(110)) xor (A(107) and B(109)) xor (A(108) and B(108)) xor (A(109) and B(107)) xor (A(110) and B(106)) xor (A(111) and B(105)) xor (A(112) and B(104)) xor (A(113) and B(103)) xor (A(114) and B(102)) xor (A(115) and B(101)) xor (A(116) and B(100)) xor (A(117) and B(99)) xor (A(118) and B(98)) xor (A(119) and B(97)) xor (A(120) and B(96)) xor (A(121) and B(95)) xor (A(122) and B(94)) xor (A(123) and B(93)) xor (A(124) and B(92)) xor (A(125) and B(91)) xor (A(126) and B(90)) xor (A(90) and B(127)) xor (A(91) and B(126)) xor (A(92) and B(125)) xor (A(93) and B(124)) xor (A(94) and B(123)) xor (A(95) and B(122)) xor (A(96) and B(121)) xor (A(97) and B(120)) xor (A(98) and B(119)) xor (A(99) and B(118)) xor (A(100) and B(117)) xor (A(101) and B(116)) xor (A(102) and B(115)) xor (A(103) and B(114)) xor (A(104) and B(113)) xor (A(105) and B(112)) xor (A(106) and B(111)) xor (A(107) and B(110)) xor (A(108) and B(109)) xor (A(109) and B(108)) xor (A(110) and B(107)) xor (A(111) and B(106)) xor (A(112) and B(105)) xor (A(113) and B(104)) xor (A(114) and B(103)) xor (A(115) and B(102)) xor (A(116) and B(101)) xor (A(117) and B(100)) xor (A(118) and B(99)) xor (A(119) and B(98)) xor (A(120) and B(97)) xor (A(121) and B(96)) xor (A(122) and B(95)) xor (A(123) and B(94)) xor (A(124) and B(93)) xor (A(125) and B(92)) xor (A(126) and B(91)) xor (A(91) and B(127)) xor (A(92) and B(126)) xor (A(93) and B(125)) xor (A(94) and B(124)) xor (A(95) and B(123)) xor (A(96) and B(122)) xor (A(97) and B(121)) xor (A(98) and B(120)) xor (A(99) and B(119)) xor (A(100) and B(118)) xor (A(101) and B(117)) xor (A(102) and B(116)) xor (A(103) and B(115)) xor (A(104) and B(114)) xor (A(105) and B(113)) xor (A(106) and B(112)) xor (A(107) and B(111)) xor (A(108) and B(110)) xor (A(109) and B(109)) xor (A(110) and B(108)) xor (A(111) and B(107)) xor (A(112) and B(106)) xor (A(113) and B(105)) xor (A(114) and B(104)) xor (A(115) and B(103)) xor (A(116) and B(102)) xor (A(117) and B(101)) xor (A(118) and B(100)) xor (A(119) and B(99)) xor (A(120) and B(98)) xor (A(121) and B(97)) xor (A(122) and B(96)) xor (A(123) and B(95)) xor (A(124) and B(94)) xor (A(125) and B(93)) xor (A(126) and B(93));
    C(92)  <= (A(0) and B(92)) xor (A(1) and B(91)) xor (A(2) and B(90)) xor (A(3) and B(89)) xor (A(4) and B(88)) xor (A(5) and B(87)) xor (A(6) and B(86)) xor (A(7) and B(85)) xor (A(8) and B(84)) xor (A(9) and B(83)) xor (A(10) and B(82)) xor (A(11) and B(81)) xor (A(12) and B(80)) xor (A(13) and B(79)) xor (A(14) and B(78)) xor (A(15) and B(77)) xor (A(16) and B(76)) xor (A(17) and B(75)) xor (A(18) and B(74)) xor (A(19) and B(73)) xor (A(20) and B(72)) xor (A(21) and B(71)) xor (A(23) and B(70)) xor (A(23) and B(69)) xor (A(24) and B(68)) xor (A(25) and B(67)) xor (A(26) and B(66)) xor (A(27) and B(65)) xor (A(28) and B(64)) xor (A(29) and B(63)) xor (A(30) and B(62)) xor (A(31) and B(61)) xor (A(32) and B(60)) xor (A(33) and B(59)) xor (A(34) and B(58)) xor (A(35) and B(57)) xor (A(36) and B(56)) xor (A(37) and B(55)) xor (A(38) and B(54)) xor (A(39) and B(53)) xor (A(40) and B(52)) xor (A(41) and B(51)) xor (A(42) and B(50)) xor (A(43) and B(49)) xor (A(44) and B(48)) xor (A(45) and B(47)) xor (A(46) and B(46)) xor (A(47) and B(45)) xor (A(48) and B(44)) xor (A(49) and B(43)) xor (A(50) and B(42)) xor (A(51) and B(41)) xor (A(52) and B(40)) xor (A(53) and B(39)) xor (A(54) and B(38)) xor (A(55) and B(37)) xor (A(56) and B(36)) xor (A(57) and B(35)) xor (A(58) and B(34)) xor (A(59) and B(33)) xor (A(60) and B(32)) xor (A(61) and B(31)) xor (A(62) and B(30)) xor (A(63) and B(29)) xor (A(64) and B(28)) xor (A(65) and B(27)) xor (A(66) and B(26)) xor (A(67) and B(25)) xor (A(68) and B(24)) xor (A(69) and B(23)) xor (A(70) and B(23)) xor (A(71) and B(21)) xor (A(72) and B(20)) xor (A(73) and B(19)) xor (A(74) and B(18)) xor (A(75) and B(17)) xor (A(76) and B(16)) xor (A(77) and B(15)) xor (A(78) and B(14)) xor (A(79) and B(13)) xor (A(80) and B(12)) xor (A(81) and B(11)) xor (A(82) and B(10)) xor (A(83) and B(9)) xor (A(84) and B(8)) xor (A(85) and B(7)) xor (A(86) and B(6)) xor (A(87) and B(5)) xor (A(88) and B(4)) xor (A(89) and B(3)) xor (A(90) and B(2)) xor (A(91) and B(1)) xor (A(92) and B(0)) xor (A(85) and B(127)) xor (A(86) and B(126)) xor (A(87) and B(125)) xor (A(88) and B(124)) xor (A(89) and B(123)) xor (A(90) and B(122)) xor (A(91) and B(121)) xor (A(92) and B(120)) xor (A(93) and B(119)) xor (A(94) and B(118)) xor (A(95) and B(117)) xor (A(96) and B(116)) xor (A(97) and B(115)) xor (A(98) and B(114)) xor (A(99) and B(113)) xor (A(100) and B(112)) xor (A(101) and B(111)) xor (A(102) and B(110)) xor (A(103) and B(109)) xor (A(104) and B(108)) xor (A(105) and B(107)) xor (A(106) and B(106)) xor (A(107) and B(105)) xor (A(108) and B(104)) xor (A(109) and B(103)) xor (A(110) and B(102)) xor (A(111) and B(101)) xor (A(112) and B(100)) xor (A(113) and B(99)) xor (A(114) and B(98)) xor (A(115) and B(97)) xor (A(116) and B(96)) xor (A(117) and B(95)) xor (A(118) and B(94)) xor (A(119) and B(93)) xor (A(120) and B(92)) xor (A(121) and B(91)) xor (A(122) and B(90)) xor (A(123) and B(89)) xor (A(124) and B(88)) xor (A(125) and B(87)) xor (A(126) and B(86)) xor (A(90) and B(127)) xor (A(91) and B(126)) xor (A(92) and B(125)) xor (A(93) and B(124)) xor (A(94) and B(123)) xor (A(95) and B(122)) xor (A(96) and B(121)) xor (A(97) and B(120)) xor (A(98) and B(119)) xor (A(99) and B(118)) xor (A(100) and B(117)) xor (A(101) and B(116)) xor (A(102) and B(115)) xor (A(103) and B(114)) xor (A(104) and B(113)) xor (A(105) and B(112)) xor (A(106) and B(111)) xor (A(107) and B(110)) xor (A(108) and B(109)) xor (A(109) and B(108)) xor (A(110) and B(107)) xor (A(111) and B(106)) xor (A(112) and B(105)) xor (A(113) and B(104)) xor (A(114) and B(103)) xor (A(115) and B(102)) xor (A(116) and B(101)) xor (A(117) and B(100)) xor (A(118) and B(99)) xor (A(119) and B(98)) xor (A(120) and B(97)) xor (A(121) and B(96)) xor (A(122) and B(95)) xor (A(123) and B(94)) xor (A(124) and B(93)) xor (A(125) and B(92)) xor (A(126) and B(91)) xor (A(91) and B(127)) xor (A(92) and B(126)) xor (A(93) and B(125)) xor (A(94) and B(124)) xor (A(95) and B(123)) xor (A(96) and B(122)) xor (A(97) and B(121)) xor (A(98) and B(120)) xor (A(99) and B(119)) xor (A(100) and B(118)) xor (A(101) and B(117)) xor (A(102) and B(116)) xor (A(103) and B(115)) xor (A(104) and B(114)) xor (A(105) and B(113)) xor (A(106) and B(112)) xor (A(107) and B(111)) xor (A(108) and B(110)) xor (A(109) and B(109)) xor (A(110) and B(108)) xor (A(111) and B(107)) xor (A(112) and B(106)) xor (A(113) and B(105)) xor (A(114) and B(104)) xor (A(115) and B(103)) xor (A(116) and B(102)) xor (A(117) and B(101)) xor (A(118) and B(100)) xor (A(119) and B(99)) xor (A(120) and B(98)) xor (A(121) and B(97)) xor (A(122) and B(96)) xor (A(123) and B(95)) xor (A(124) and B(94)) xor (A(125) and B(93)) xor (A(126) and B(92)) xor (A(92) and B(127)) xor (A(93) and B(126)) xor (A(94) and B(125)) xor (A(95) and B(124)) xor (A(96) and B(123)) xor (A(97) and B(122)) xor (A(98) and B(121)) xor (A(99) and B(120)) xor (A(100) and B(119)) xor (A(101) and B(118)) xor (A(102) and B(117)) xor (A(103) and B(116)) xor (A(104) and B(115)) xor (A(105) and B(114)) xor (A(106) and B(113)) xor (A(107) and B(112)) xor (A(108) and B(111)) xor (A(109) and B(110)) xor (A(110) and B(109)) xor (A(111) and B(108)) xor (A(112) and B(107)) xor (A(113) and B(106)) xor (A(114) and B(105)) xor (A(115) and B(104)) xor (A(116) and B(103)) xor (A(117) and B(102)) xor (A(118) and B(101)) xor (A(119) and B(100)) xor (A(120) and B(99)) xor (A(121) and B(98)) xor (A(122) and B(97)) xor (A(123) and B(96)) xor (A(124) and B(95)) xor (A(125) and B(94)) xor (A(126) and B(94));
    C(93)  <= (A(0) and B(93)) xor (A(1) and B(92)) xor (A(2) and B(91)) xor (A(3) and B(90)) xor (A(4) and B(89)) xor (A(5) and B(88)) xor (A(6) and B(87)) xor (A(7) and B(86)) xor (A(8) and B(85)) xor (A(9) and B(84)) xor (A(10) and B(83)) xor (A(11) and B(82)) xor (A(12) and B(81)) xor (A(13) and B(80)) xor (A(14) and B(79)) xor (A(15) and B(78)) xor (A(16) and B(77)) xor (A(17) and B(76)) xor (A(18) and B(75)) xor (A(19) and B(74)) xor (A(20) and B(73)) xor (A(21) and B(72)) xor (A(23) and B(71)) xor (A(23) and B(70)) xor (A(24) and B(69)) xor (A(25) and B(68)) xor (A(26) and B(67)) xor (A(27) and B(66)) xor (A(28) and B(65)) xor (A(29) and B(64)) xor (A(30) and B(63)) xor (A(31) and B(62)) xor (A(32) and B(61)) xor (A(33) and B(60)) xor (A(34) and B(59)) xor (A(35) and B(58)) xor (A(36) and B(57)) xor (A(37) and B(56)) xor (A(38) and B(55)) xor (A(39) and B(54)) xor (A(40) and B(53)) xor (A(41) and B(52)) xor (A(42) and B(51)) xor (A(43) and B(50)) xor (A(44) and B(49)) xor (A(45) and B(48)) xor (A(46) and B(47)) xor (A(47) and B(46)) xor (A(48) and B(45)) xor (A(49) and B(44)) xor (A(50) and B(43)) xor (A(51) and B(42)) xor (A(52) and B(41)) xor (A(53) and B(40)) xor (A(54) and B(39)) xor (A(55) and B(38)) xor (A(56) and B(37)) xor (A(57) and B(36)) xor (A(58) and B(35)) xor (A(59) and B(34)) xor (A(60) and B(33)) xor (A(61) and B(32)) xor (A(62) and B(31)) xor (A(63) and B(30)) xor (A(64) and B(29)) xor (A(65) and B(28)) xor (A(66) and B(27)) xor (A(67) and B(26)) xor (A(68) and B(25)) xor (A(69) and B(24)) xor (A(70) and B(23)) xor (A(71) and B(23)) xor (A(72) and B(21)) xor (A(73) and B(20)) xor (A(74) and B(19)) xor (A(75) and B(18)) xor (A(76) and B(17)) xor (A(77) and B(16)) xor (A(78) and B(15)) xor (A(79) and B(14)) xor (A(80) and B(13)) xor (A(81) and B(12)) xor (A(82) and B(11)) xor (A(83) and B(10)) xor (A(84) and B(9)) xor (A(85) and B(8)) xor (A(86) and B(7)) xor (A(87) and B(6)) xor (A(88) and B(5)) xor (A(89) and B(4)) xor (A(90) and B(3)) xor (A(91) and B(2)) xor (A(92) and B(1)) xor (A(93) and B(0)) xor (A(86) and B(127)) xor (A(87) and B(126)) xor (A(88) and B(125)) xor (A(89) and B(124)) xor (A(90) and B(123)) xor (A(91) and B(122)) xor (A(92) and B(121)) xor (A(93) and B(120)) xor (A(94) and B(119)) xor (A(95) and B(118)) xor (A(96) and B(117)) xor (A(97) and B(116)) xor (A(98) and B(115)) xor (A(99) and B(114)) xor (A(100) and B(113)) xor (A(101) and B(112)) xor (A(102) and B(111)) xor (A(103) and B(110)) xor (A(104) and B(109)) xor (A(105) and B(108)) xor (A(106) and B(107)) xor (A(107) and B(106)) xor (A(108) and B(105)) xor (A(109) and B(104)) xor (A(110) and B(103)) xor (A(111) and B(102)) xor (A(112) and B(101)) xor (A(113) and B(100)) xor (A(114) and B(99)) xor (A(115) and B(98)) xor (A(116) and B(97)) xor (A(117) and B(96)) xor (A(118) and B(95)) xor (A(119) and B(94)) xor (A(120) and B(93)) xor (A(121) and B(92)) xor (A(122) and B(91)) xor (A(123) and B(90)) xor (A(124) and B(89)) xor (A(125) and B(88)) xor (A(126) and B(87)) xor (A(91) and B(127)) xor (A(92) and B(126)) xor (A(93) and B(125)) xor (A(94) and B(124)) xor (A(95) and B(123)) xor (A(96) and B(122)) xor (A(97) and B(121)) xor (A(98) and B(120)) xor (A(99) and B(119)) xor (A(100) and B(118)) xor (A(101) and B(117)) xor (A(102) and B(116)) xor (A(103) and B(115)) xor (A(104) and B(114)) xor (A(105) and B(113)) xor (A(106) and B(112)) xor (A(107) and B(111)) xor (A(108) and B(110)) xor (A(109) and B(109)) xor (A(110) and B(108)) xor (A(111) and B(107)) xor (A(112) and B(106)) xor (A(113) and B(105)) xor (A(114) and B(104)) xor (A(115) and B(103)) xor (A(116) and B(102)) xor (A(117) and B(101)) xor (A(118) and B(100)) xor (A(119) and B(99)) xor (A(120) and B(98)) xor (A(121) and B(97)) xor (A(122) and B(96)) xor (A(123) and B(95)) xor (A(124) and B(94)) xor (A(125) and B(93)) xor (A(126) and B(92)) xor (A(92) and B(127)) xor (A(93) and B(126)) xor (A(94) and B(125)) xor (A(95) and B(124)) xor (A(96) and B(123)) xor (A(97) and B(122)) xor (A(98) and B(121)) xor (A(99) and B(120)) xor (A(100) and B(119)) xor (A(101) and B(118)) xor (A(102) and B(117)) xor (A(103) and B(116)) xor (A(104) and B(115)) xor (A(105) and B(114)) xor (A(106) and B(113)) xor (A(107) and B(112)) xor (A(108) and B(111)) xor (A(109) and B(110)) xor (A(110) and B(109)) xor (A(111) and B(108)) xor (A(112) and B(107)) xor (A(113) and B(106)) xor (A(114) and B(105)) xor (A(115) and B(104)) xor (A(116) and B(103)) xor (A(117) and B(102)) xor (A(118) and B(101)) xor (A(119) and B(100)) xor (A(120) and B(99)) xor (A(121) and B(98)) xor (A(122) and B(97)) xor (A(123) and B(96)) xor (A(124) and B(95)) xor (A(125) and B(94)) xor (A(126) and B(93)) xor (A(93) and B(127)) xor (A(94) and B(126)) xor (A(95) and B(125)) xor (A(96) and B(124)) xor (A(97) and B(123)) xor (A(98) and B(122)) xor (A(99) and B(121)) xor (A(100) and B(120)) xor (A(101) and B(119)) xor (A(102) and B(118)) xor (A(103) and B(117)) xor (A(104) and B(116)) xor (A(105) and B(115)) xor (A(106) and B(114)) xor (A(107) and B(113)) xor (A(108) and B(112)) xor (A(109) and B(111)) xor (A(110) and B(110)) xor (A(111) and B(109)) xor (A(112) and B(108)) xor (A(113) and B(107)) xor (A(114) and B(106)) xor (A(115) and B(105)) xor (A(116) and B(104)) xor (A(117) and B(103)) xor (A(118) and B(102)) xor (A(119) and B(101)) xor (A(120) and B(100)) xor (A(121) and B(99)) xor (A(122) and B(98)) xor (A(123) and B(97)) xor (A(124) and B(96)) xor (A(125) and B(95)) xor (A(126) and B(95));
    C(94)  <= (A(0) and B(94)) xor (A(1) and B(93)) xor (A(2) and B(92)) xor (A(3) and B(91)) xor (A(4) and B(90)) xor (A(5) and B(89)) xor (A(6) and B(88)) xor (A(7) and B(87)) xor (A(8) and B(86)) xor (A(9) and B(85)) xor (A(10) and B(84)) xor (A(11) and B(83)) xor (A(12) and B(82)) xor (A(13) and B(81)) xor (A(14) and B(80)) xor (A(15) and B(79)) xor (A(16) and B(78)) xor (A(17) and B(77)) xor (A(18) and B(76)) xor (A(19) and B(75)) xor (A(20) and B(74)) xor (A(21) and B(73)) xor (A(23) and B(72)) xor (A(23) and B(71)) xor (A(24) and B(70)) xor (A(25) and B(69)) xor (A(26) and B(68)) xor (A(27) and B(67)) xor (A(28) and B(66)) xor (A(29) and B(65)) xor (A(30) and B(64)) xor (A(31) and B(63)) xor (A(32) and B(62)) xor (A(33) and B(61)) xor (A(34) and B(60)) xor (A(35) and B(59)) xor (A(36) and B(58)) xor (A(37) and B(57)) xor (A(38) and B(56)) xor (A(39) and B(55)) xor (A(40) and B(54)) xor (A(41) and B(53)) xor (A(42) and B(52)) xor (A(43) and B(51)) xor (A(44) and B(50)) xor (A(45) and B(49)) xor (A(46) and B(48)) xor (A(47) and B(47)) xor (A(48) and B(46)) xor (A(49) and B(45)) xor (A(50) and B(44)) xor (A(51) and B(43)) xor (A(52) and B(42)) xor (A(53) and B(41)) xor (A(54) and B(40)) xor (A(55) and B(39)) xor (A(56) and B(38)) xor (A(57) and B(37)) xor (A(58) and B(36)) xor (A(59) and B(35)) xor (A(60) and B(34)) xor (A(61) and B(33)) xor (A(62) and B(32)) xor (A(63) and B(31)) xor (A(64) and B(30)) xor (A(65) and B(29)) xor (A(66) and B(28)) xor (A(67) and B(27)) xor (A(68) and B(26)) xor (A(69) and B(25)) xor (A(70) and B(24)) xor (A(71) and B(23)) xor (A(72) and B(23)) xor (A(73) and B(21)) xor (A(74) and B(20)) xor (A(75) and B(19)) xor (A(76) and B(18)) xor (A(77) and B(17)) xor (A(78) and B(16)) xor (A(79) and B(15)) xor (A(80) and B(14)) xor (A(81) and B(13)) xor (A(82) and B(12)) xor (A(83) and B(11)) xor (A(84) and B(10)) xor (A(85) and B(9)) xor (A(86) and B(8)) xor (A(87) and B(7)) xor (A(88) and B(6)) xor (A(89) and B(5)) xor (A(90) and B(4)) xor (A(91) and B(3)) xor (A(92) and B(2)) xor (A(93) and B(1)) xor (A(94) and B(0)) xor (A(87) and B(127)) xor (A(88) and B(126)) xor (A(89) and B(125)) xor (A(90) and B(124)) xor (A(91) and B(123)) xor (A(92) and B(122)) xor (A(93) and B(121)) xor (A(94) and B(120)) xor (A(95) and B(119)) xor (A(96) and B(118)) xor (A(97) and B(117)) xor (A(98) and B(116)) xor (A(99) and B(115)) xor (A(100) and B(114)) xor (A(101) and B(113)) xor (A(102) and B(112)) xor (A(103) and B(111)) xor (A(104) and B(110)) xor (A(105) and B(109)) xor (A(106) and B(108)) xor (A(107) and B(107)) xor (A(108) and B(106)) xor (A(109) and B(105)) xor (A(110) and B(104)) xor (A(111) and B(103)) xor (A(112) and B(102)) xor (A(113) and B(101)) xor (A(114) and B(100)) xor (A(115) and B(99)) xor (A(116) and B(98)) xor (A(117) and B(97)) xor (A(118) and B(96)) xor (A(119) and B(95)) xor (A(120) and B(94)) xor (A(121) and B(93)) xor (A(122) and B(92)) xor (A(123) and B(91)) xor (A(124) and B(90)) xor (A(125) and B(89)) xor (A(126) and B(88)) xor (A(92) and B(127)) xor (A(93) and B(126)) xor (A(94) and B(125)) xor (A(95) and B(124)) xor (A(96) and B(123)) xor (A(97) and B(122)) xor (A(98) and B(121)) xor (A(99) and B(120)) xor (A(100) and B(119)) xor (A(101) and B(118)) xor (A(102) and B(117)) xor (A(103) and B(116)) xor (A(104) and B(115)) xor (A(105) and B(114)) xor (A(106) and B(113)) xor (A(107) and B(112)) xor (A(108) and B(111)) xor (A(109) and B(110)) xor (A(110) and B(109)) xor (A(111) and B(108)) xor (A(112) and B(107)) xor (A(113) and B(106)) xor (A(114) and B(105)) xor (A(115) and B(104)) xor (A(116) and B(103)) xor (A(117) and B(102)) xor (A(118) and B(101)) xor (A(119) and B(100)) xor (A(120) and B(99)) xor (A(121) and B(98)) xor (A(122) and B(97)) xor (A(123) and B(96)) xor (A(124) and B(95)) xor (A(125) and B(94)) xor (A(126) and B(93)) xor (A(93) and B(127)) xor (A(94) and B(126)) xor (A(95) and B(125)) xor (A(96) and B(124)) xor (A(97) and B(123)) xor (A(98) and B(122)) xor (A(99) and B(121)) xor (A(100) and B(120)) xor (A(101) and B(119)) xor (A(102) and B(118)) xor (A(103) and B(117)) xor (A(104) and B(116)) xor (A(105) and B(115)) xor (A(106) and B(114)) xor (A(107) and B(113)) xor (A(108) and B(112)) xor (A(109) and B(111)) xor (A(110) and B(110)) xor (A(111) and B(109)) xor (A(112) and B(108)) xor (A(113) and B(107)) xor (A(114) and B(106)) xor (A(115) and B(105)) xor (A(116) and B(104)) xor (A(117) and B(103)) xor (A(118) and B(102)) xor (A(119) and B(101)) xor (A(120) and B(100)) xor (A(121) and B(99)) xor (A(122) and B(98)) xor (A(123) and B(97)) xor (A(124) and B(96)) xor (A(125) and B(95)) xor (A(126) and B(94)) xor (A(94) and B(127)) xor (A(95) and B(126)) xor (A(96) and B(125)) xor (A(97) and B(124)) xor (A(98) and B(123)) xor (A(99) and B(122)) xor (A(100) and B(121)) xor (A(101) and B(120)) xor (A(102) and B(119)) xor (A(103) and B(118)) xor (A(104) and B(117)) xor (A(105) and B(116)) xor (A(106) and B(115)) xor (A(107) and B(114)) xor (A(108) and B(113)) xor (A(109) and B(112)) xor (A(110) and B(111)) xor (A(111) and B(110)) xor (A(112) and B(109)) xor (A(113) and B(108)) xor (A(114) and B(107)) xor (A(115) and B(106)) xor (A(116) and B(105)) xor (A(117) and B(104)) xor (A(118) and B(103)) xor (A(119) and B(102)) xor (A(120) and B(101)) xor (A(121) and B(100)) xor (A(122) and B(99)) xor (A(123) and B(98)) xor (A(124) and B(97)) xor (A(125) and B(96)) xor (A(126) and B(96));
    C(95)  <= (A(0) and B(95)) xor (A(1) and B(94)) xor (A(2) and B(93)) xor (A(3) and B(92)) xor (A(4) and B(91)) xor (A(5) and B(90)) xor (A(6) and B(89)) xor (A(7) and B(88)) xor (A(8) and B(87)) xor (A(9) and B(86)) xor (A(10) and B(85)) xor (A(11) and B(84)) xor (A(12) and B(83)) xor (A(13) and B(82)) xor (A(14) and B(81)) xor (A(15) and B(80)) xor (A(16) and B(79)) xor (A(17) and B(78)) xor (A(18) and B(77)) xor (A(19) and B(76)) xor (A(20) and B(75)) xor (A(21) and B(74)) xor (A(23) and B(73)) xor (A(23) and B(72)) xor (A(24) and B(71)) xor (A(25) and B(70)) xor (A(26) and B(69)) xor (A(27) and B(68)) xor (A(28) and B(67)) xor (A(29) and B(66)) xor (A(30) and B(65)) xor (A(31) and B(64)) xor (A(32) and B(63)) xor (A(33) and B(62)) xor (A(34) and B(61)) xor (A(35) and B(60)) xor (A(36) and B(59)) xor (A(37) and B(58)) xor (A(38) and B(57)) xor (A(39) and B(56)) xor (A(40) and B(55)) xor (A(41) and B(54)) xor (A(42) and B(53)) xor (A(43) and B(52)) xor (A(44) and B(51)) xor (A(45) and B(50)) xor (A(46) and B(49)) xor (A(47) and B(48)) xor (A(48) and B(47)) xor (A(49) and B(46)) xor (A(50) and B(45)) xor (A(51) and B(44)) xor (A(52) and B(43)) xor (A(53) and B(42)) xor (A(54) and B(41)) xor (A(55) and B(40)) xor (A(56) and B(39)) xor (A(57) and B(38)) xor (A(58) and B(37)) xor (A(59) and B(36)) xor (A(60) and B(35)) xor (A(61) and B(34)) xor (A(62) and B(33)) xor (A(63) and B(32)) xor (A(64) and B(31)) xor (A(65) and B(30)) xor (A(66) and B(29)) xor (A(67) and B(28)) xor (A(68) and B(27)) xor (A(69) and B(26)) xor (A(70) and B(25)) xor (A(71) and B(24)) xor (A(72) and B(23)) xor (A(73) and B(23)) xor (A(74) and B(21)) xor (A(75) and B(20)) xor (A(76) and B(19)) xor (A(77) and B(18)) xor (A(78) and B(17)) xor (A(79) and B(16)) xor (A(80) and B(15)) xor (A(81) and B(14)) xor (A(82) and B(13)) xor (A(83) and B(12)) xor (A(84) and B(11)) xor (A(85) and B(10)) xor (A(86) and B(9)) xor (A(87) and B(8)) xor (A(88) and B(7)) xor (A(89) and B(6)) xor (A(90) and B(5)) xor (A(91) and B(4)) xor (A(92) and B(3)) xor (A(93) and B(2)) xor (A(94) and B(1)) xor (A(95) and B(0)) xor (A(88) and B(127)) xor (A(89) and B(126)) xor (A(90) and B(125)) xor (A(91) and B(124)) xor (A(92) and B(123)) xor (A(93) and B(122)) xor (A(94) and B(121)) xor (A(95) and B(120)) xor (A(96) and B(119)) xor (A(97) and B(118)) xor (A(98) and B(117)) xor (A(99) and B(116)) xor (A(100) and B(115)) xor (A(101) and B(114)) xor (A(102) and B(113)) xor (A(103) and B(112)) xor (A(104) and B(111)) xor (A(105) and B(110)) xor (A(106) and B(109)) xor (A(107) and B(108)) xor (A(108) and B(107)) xor (A(109) and B(106)) xor (A(110) and B(105)) xor (A(111) and B(104)) xor (A(112) and B(103)) xor (A(113) and B(102)) xor (A(114) and B(101)) xor (A(115) and B(100)) xor (A(116) and B(99)) xor (A(117) and B(98)) xor (A(118) and B(97)) xor (A(119) and B(96)) xor (A(120) and B(95)) xor (A(121) and B(94)) xor (A(122) and B(93)) xor (A(123) and B(92)) xor (A(124) and B(91)) xor (A(125) and B(90)) xor (A(126) and B(89)) xor (A(93) and B(127)) xor (A(94) and B(126)) xor (A(95) and B(125)) xor (A(96) and B(124)) xor (A(97) and B(123)) xor (A(98) and B(122)) xor (A(99) and B(121)) xor (A(100) and B(120)) xor (A(101) and B(119)) xor (A(102) and B(118)) xor (A(103) and B(117)) xor (A(104) and B(116)) xor (A(105) and B(115)) xor (A(106) and B(114)) xor (A(107) and B(113)) xor (A(108) and B(112)) xor (A(109) and B(111)) xor (A(110) and B(110)) xor (A(111) and B(109)) xor (A(112) and B(108)) xor (A(113) and B(107)) xor (A(114) and B(106)) xor (A(115) and B(105)) xor (A(116) and B(104)) xor (A(117) and B(103)) xor (A(118) and B(102)) xor (A(119) and B(101)) xor (A(120) and B(100)) xor (A(121) and B(99)) xor (A(122) and B(98)) xor (A(123) and B(97)) xor (A(124) and B(96)) xor (A(125) and B(95)) xor (A(126) and B(94)) xor (A(94) and B(127)) xor (A(95) and B(126)) xor (A(96) and B(125)) xor (A(97) and B(124)) xor (A(98) and B(123)) xor (A(99) and B(122)) xor (A(100) and B(121)) xor (A(101) and B(120)) xor (A(102) and B(119)) xor (A(103) and B(118)) xor (A(104) and B(117)) xor (A(105) and B(116)) xor (A(106) and B(115)) xor (A(107) and B(114)) xor (A(108) and B(113)) xor (A(109) and B(112)) xor (A(110) and B(111)) xor (A(111) and B(110)) xor (A(112) and B(109)) xor (A(113) and B(108)) xor (A(114) and B(107)) xor (A(115) and B(106)) xor (A(116) and B(105)) xor (A(117) and B(104)) xor (A(118) and B(103)) xor (A(119) and B(102)) xor (A(120) and B(101)) xor (A(121) and B(100)) xor (A(122) and B(99)) xor (A(123) and B(98)) xor (A(124) and B(97)) xor (A(125) and B(96)) xor (A(126) and B(95)) xor (A(95) and B(127)) xor (A(96) and B(126)) xor (A(97) and B(125)) xor (A(98) and B(124)) xor (A(99) and B(123)) xor (A(100) and B(122)) xor (A(101) and B(121)) xor (A(102) and B(120)) xor (A(103) and B(119)) xor (A(104) and B(118)) xor (A(105) and B(117)) xor (A(106) and B(116)) xor (A(107) and B(115)) xor (A(108) and B(114)) xor (A(109) and B(113)) xor (A(110) and B(112)) xor (A(111) and B(111)) xor (A(112) and B(110)) xor (A(113) and B(109)) xor (A(114) and B(108)) xor (A(115) and B(107)) xor (A(116) and B(106)) xor (A(117) and B(105)) xor (A(118) and B(104)) xor (A(119) and B(103)) xor (A(120) and B(102)) xor (A(121) and B(101)) xor (A(122) and B(100)) xor (A(123) and B(99)) xor (A(124) and B(98)) xor (A(125) and B(97)) xor (A(126) and B(97));
    C(96)  <= (A(0) and B(96)) xor (A(1) and B(95)) xor (A(2) and B(94)) xor (A(3) and B(93)) xor (A(4) and B(92)) xor (A(5) and B(91)) xor (A(6) and B(90)) xor (A(7) and B(89)) xor (A(8) and B(88)) xor (A(9) and B(87)) xor (A(10) and B(86)) xor (A(11) and B(85)) xor (A(12) and B(84)) xor (A(13) and B(83)) xor (A(14) and B(82)) xor (A(15) and B(81)) xor (A(16) and B(80)) xor (A(17) and B(79)) xor (A(18) and B(78)) xor (A(19) and B(77)) xor (A(20) and B(76)) xor (A(21) and B(75)) xor (A(23) and B(74)) xor (A(23) and B(73)) xor (A(24) and B(72)) xor (A(25) and B(71)) xor (A(26) and B(70)) xor (A(27) and B(69)) xor (A(28) and B(68)) xor (A(29) and B(67)) xor (A(30) and B(66)) xor (A(31) and B(65)) xor (A(32) and B(64)) xor (A(33) and B(63)) xor (A(34) and B(62)) xor (A(35) and B(61)) xor (A(36) and B(60)) xor (A(37) and B(59)) xor (A(38) and B(58)) xor (A(39) and B(57)) xor (A(40) and B(56)) xor (A(41) and B(55)) xor (A(42) and B(54)) xor (A(43) and B(53)) xor (A(44) and B(52)) xor (A(45) and B(51)) xor (A(46) and B(50)) xor (A(47) and B(49)) xor (A(48) and B(48)) xor (A(49) and B(47)) xor (A(50) and B(46)) xor (A(51) and B(45)) xor (A(52) and B(44)) xor (A(53) and B(43)) xor (A(54) and B(42)) xor (A(55) and B(41)) xor (A(56) and B(40)) xor (A(57) and B(39)) xor (A(58) and B(38)) xor (A(59) and B(37)) xor (A(60) and B(36)) xor (A(61) and B(35)) xor (A(62) and B(34)) xor (A(63) and B(33)) xor (A(64) and B(32)) xor (A(65) and B(31)) xor (A(66) and B(30)) xor (A(67) and B(29)) xor (A(68) and B(28)) xor (A(69) and B(27)) xor (A(70) and B(26)) xor (A(71) and B(25)) xor (A(72) and B(24)) xor (A(73) and B(23)) xor (A(74) and B(23)) xor (A(75) and B(21)) xor (A(76) and B(20)) xor (A(77) and B(19)) xor (A(78) and B(18)) xor (A(79) and B(17)) xor (A(80) and B(16)) xor (A(81) and B(15)) xor (A(82) and B(14)) xor (A(83) and B(13)) xor (A(84) and B(12)) xor (A(85) and B(11)) xor (A(86) and B(10)) xor (A(87) and B(9)) xor (A(88) and B(8)) xor (A(89) and B(7)) xor (A(90) and B(6)) xor (A(91) and B(5)) xor (A(92) and B(4)) xor (A(93) and B(3)) xor (A(94) and B(2)) xor (A(95) and B(1)) xor (A(96) and B(0)) xor (A(89) and B(127)) xor (A(90) and B(126)) xor (A(91) and B(125)) xor (A(92) and B(124)) xor (A(93) and B(123)) xor (A(94) and B(122)) xor (A(95) and B(121)) xor (A(96) and B(120)) xor (A(97) and B(119)) xor (A(98) and B(118)) xor (A(99) and B(117)) xor (A(100) and B(116)) xor (A(101) and B(115)) xor (A(102) and B(114)) xor (A(103) and B(113)) xor (A(104) and B(112)) xor (A(105) and B(111)) xor (A(106) and B(110)) xor (A(107) and B(109)) xor (A(108) and B(108)) xor (A(109) and B(107)) xor (A(110) and B(106)) xor (A(111) and B(105)) xor (A(112) and B(104)) xor (A(113) and B(103)) xor (A(114) and B(102)) xor (A(115) and B(101)) xor (A(116) and B(100)) xor (A(117) and B(99)) xor (A(118) and B(98)) xor (A(119) and B(97)) xor (A(120) and B(96)) xor (A(121) and B(95)) xor (A(122) and B(94)) xor (A(123) and B(93)) xor (A(124) and B(92)) xor (A(125) and B(91)) xor (A(126) and B(90)) xor (A(94) and B(127)) xor (A(95) and B(126)) xor (A(96) and B(125)) xor (A(97) and B(124)) xor (A(98) and B(123)) xor (A(99) and B(122)) xor (A(100) and B(121)) xor (A(101) and B(120)) xor (A(102) and B(119)) xor (A(103) and B(118)) xor (A(104) and B(117)) xor (A(105) and B(116)) xor (A(106) and B(115)) xor (A(107) and B(114)) xor (A(108) and B(113)) xor (A(109) and B(112)) xor (A(110) and B(111)) xor (A(111) and B(110)) xor (A(112) and B(109)) xor (A(113) and B(108)) xor (A(114) and B(107)) xor (A(115) and B(106)) xor (A(116) and B(105)) xor (A(117) and B(104)) xor (A(118) and B(103)) xor (A(119) and B(102)) xor (A(120) and B(101)) xor (A(121) and B(100)) xor (A(122) and B(99)) xor (A(123) and B(98)) xor (A(124) and B(97)) xor (A(125) and B(96)) xor (A(126) and B(95)) xor (A(95) and B(127)) xor (A(96) and B(126)) xor (A(97) and B(125)) xor (A(98) and B(124)) xor (A(99) and B(123)) xor (A(100) and B(122)) xor (A(101) and B(121)) xor (A(102) and B(120)) xor (A(103) and B(119)) xor (A(104) and B(118)) xor (A(105) and B(117)) xor (A(106) and B(116)) xor (A(107) and B(115)) xor (A(108) and B(114)) xor (A(109) and B(113)) xor (A(110) and B(112)) xor (A(111) and B(111)) xor (A(112) and B(110)) xor (A(113) and B(109)) xor (A(114) and B(108)) xor (A(115) and B(107)) xor (A(116) and B(106)) xor (A(117) and B(105)) xor (A(118) and B(104)) xor (A(119) and B(103)) xor (A(120) and B(102)) xor (A(121) and B(101)) xor (A(122) and B(100)) xor (A(123) and B(99)) xor (A(124) and B(98)) xor (A(125) and B(97)) xor (A(126) and B(96)) xor (A(96) and B(127)) xor (A(97) and B(126)) xor (A(98) and B(125)) xor (A(99) and B(124)) xor (A(100) and B(123)) xor (A(101) and B(122)) xor (A(102) and B(121)) xor (A(103) and B(120)) xor (A(104) and B(119)) xor (A(105) and B(118)) xor (A(106) and B(117)) xor (A(107) and B(116)) xor (A(108) and B(115)) xor (A(109) and B(114)) xor (A(110) and B(113)) xor (A(111) and B(112)) xor (A(112) and B(111)) xor (A(113) and B(110)) xor (A(114) and B(109)) xor (A(115) and B(108)) xor (A(116) and B(107)) xor (A(117) and B(106)) xor (A(118) and B(105)) xor (A(119) and B(104)) xor (A(120) and B(103)) xor (A(121) and B(102)) xor (A(122) and B(101)) xor (A(123) and B(100)) xor (A(124) and B(99)) xor (A(125) and B(98)) xor (A(126) and B(98));
    C(97)  <= (A(0) and B(97)) xor (A(1) and B(96)) xor (A(2) and B(95)) xor (A(3) and B(94)) xor (A(4) and B(93)) xor (A(5) and B(92)) xor (A(6) and B(91)) xor (A(7) and B(90)) xor (A(8) and B(89)) xor (A(9) and B(88)) xor (A(10) and B(87)) xor (A(11) and B(86)) xor (A(12) and B(85)) xor (A(13) and B(84)) xor (A(14) and B(83)) xor (A(15) and B(82)) xor (A(16) and B(81)) xor (A(17) and B(80)) xor (A(18) and B(79)) xor (A(19) and B(78)) xor (A(20) and B(77)) xor (A(21) and B(76)) xor (A(23) and B(75)) xor (A(23) and B(74)) xor (A(24) and B(73)) xor (A(25) and B(72)) xor (A(26) and B(71)) xor (A(27) and B(70)) xor (A(28) and B(69)) xor (A(29) and B(68)) xor (A(30) and B(67)) xor (A(31) and B(66)) xor (A(32) and B(65)) xor (A(33) and B(64)) xor (A(34) and B(63)) xor (A(35) and B(62)) xor (A(36) and B(61)) xor (A(37) and B(60)) xor (A(38) and B(59)) xor (A(39) and B(58)) xor (A(40) and B(57)) xor (A(41) and B(56)) xor (A(42) and B(55)) xor (A(43) and B(54)) xor (A(44) and B(53)) xor (A(45) and B(52)) xor (A(46) and B(51)) xor (A(47) and B(50)) xor (A(48) and B(49)) xor (A(49) and B(48)) xor (A(50) and B(47)) xor (A(51) and B(46)) xor (A(52) and B(45)) xor (A(53) and B(44)) xor (A(54) and B(43)) xor (A(55) and B(42)) xor (A(56) and B(41)) xor (A(57) and B(40)) xor (A(58) and B(39)) xor (A(59) and B(38)) xor (A(60) and B(37)) xor (A(61) and B(36)) xor (A(62) and B(35)) xor (A(63) and B(34)) xor (A(64) and B(33)) xor (A(65) and B(32)) xor (A(66) and B(31)) xor (A(67) and B(30)) xor (A(68) and B(29)) xor (A(69) and B(28)) xor (A(70) and B(27)) xor (A(71) and B(26)) xor (A(72) and B(25)) xor (A(73) and B(24)) xor (A(74) and B(23)) xor (A(75) and B(23)) xor (A(76) and B(21)) xor (A(77) and B(20)) xor (A(78) and B(19)) xor (A(79) and B(18)) xor (A(80) and B(17)) xor (A(81) and B(16)) xor (A(82) and B(15)) xor (A(83) and B(14)) xor (A(84) and B(13)) xor (A(85) and B(12)) xor (A(86) and B(11)) xor (A(87) and B(10)) xor (A(88) and B(9)) xor (A(89) and B(8)) xor (A(90) and B(7)) xor (A(91) and B(6)) xor (A(92) and B(5)) xor (A(93) and B(4)) xor (A(94) and B(3)) xor (A(95) and B(2)) xor (A(96) and B(1)) xor (A(97) and B(0)) xor (A(90) and B(127)) xor (A(91) and B(126)) xor (A(92) and B(125)) xor (A(93) and B(124)) xor (A(94) and B(123)) xor (A(95) and B(122)) xor (A(96) and B(121)) xor (A(97) and B(120)) xor (A(98) and B(119)) xor (A(99) and B(118)) xor (A(100) and B(117)) xor (A(101) and B(116)) xor (A(102) and B(115)) xor (A(103) and B(114)) xor (A(104) and B(113)) xor (A(105) and B(112)) xor (A(106) and B(111)) xor (A(107) and B(110)) xor (A(108) and B(109)) xor (A(109) and B(108)) xor (A(110) and B(107)) xor (A(111) and B(106)) xor (A(112) and B(105)) xor (A(113) and B(104)) xor (A(114) and B(103)) xor (A(115) and B(102)) xor (A(116) and B(101)) xor (A(117) and B(100)) xor (A(118) and B(99)) xor (A(119) and B(98)) xor (A(120) and B(97)) xor (A(121) and B(96)) xor (A(122) and B(95)) xor (A(123) and B(94)) xor (A(124) and B(93)) xor (A(125) and B(92)) xor (A(126) and B(91)) xor (A(95) and B(127)) xor (A(96) and B(126)) xor (A(97) and B(125)) xor (A(98) and B(124)) xor (A(99) and B(123)) xor (A(100) and B(122)) xor (A(101) and B(121)) xor (A(102) and B(120)) xor (A(103) and B(119)) xor (A(104) and B(118)) xor (A(105) and B(117)) xor (A(106) and B(116)) xor (A(107) and B(115)) xor (A(108) and B(114)) xor (A(109) and B(113)) xor (A(110) and B(112)) xor (A(111) and B(111)) xor (A(112) and B(110)) xor (A(113) and B(109)) xor (A(114) and B(108)) xor (A(115) and B(107)) xor (A(116) and B(106)) xor (A(117) and B(105)) xor (A(118) and B(104)) xor (A(119) and B(103)) xor (A(120) and B(102)) xor (A(121) and B(101)) xor (A(122) and B(100)) xor (A(123) and B(99)) xor (A(124) and B(98)) xor (A(125) and B(97)) xor (A(126) and B(96)) xor (A(96) and B(127)) xor (A(97) and B(126)) xor (A(98) and B(125)) xor (A(99) and B(124)) xor (A(100) and B(123)) xor (A(101) and B(122)) xor (A(102) and B(121)) xor (A(103) and B(120)) xor (A(104) and B(119)) xor (A(105) and B(118)) xor (A(106) and B(117)) xor (A(107) and B(116)) xor (A(108) and B(115)) xor (A(109) and B(114)) xor (A(110) and B(113)) xor (A(111) and B(112)) xor (A(112) and B(111)) xor (A(113) and B(110)) xor (A(114) and B(109)) xor (A(115) and B(108)) xor (A(116) and B(107)) xor (A(117) and B(106)) xor (A(118) and B(105)) xor (A(119) and B(104)) xor (A(120) and B(103)) xor (A(121) and B(102)) xor (A(122) and B(101)) xor (A(123) and B(100)) xor (A(124) and B(99)) xor (A(125) and B(98)) xor (A(126) and B(97)) xor (A(97) and B(127)) xor (A(98) and B(126)) xor (A(99) and B(125)) xor (A(100) and B(124)) xor (A(101) and B(123)) xor (A(102) and B(122)) xor (A(103) and B(121)) xor (A(104) and B(120)) xor (A(105) and B(119)) xor (A(106) and B(118)) xor (A(107) and B(117)) xor (A(108) and B(116)) xor (A(109) and B(115)) xor (A(110) and B(114)) xor (A(111) and B(113)) xor (A(112) and B(112)) xor (A(113) and B(111)) xor (A(114) and B(110)) xor (A(115) and B(109)) xor (A(116) and B(108)) xor (A(117) and B(107)) xor (A(118) and B(106)) xor (A(119) and B(105)) xor (A(120) and B(104)) xor (A(121) and B(103)) xor (A(122) and B(102)) xor (A(123) and B(101)) xor (A(124) and B(100)) xor (A(125) and B(99)) xor (A(126) and B(99));
    C(98)  <= (A(0) and B(98)) xor (A(1) and B(97)) xor (A(2) and B(96)) xor (A(3) and B(95)) xor (A(4) and B(94)) xor (A(5) and B(93)) xor (A(6) and B(92)) xor (A(7) and B(91)) xor (A(8) and B(90)) xor (A(9) and B(89)) xor (A(10) and B(88)) xor (A(11) and B(87)) xor (A(12) and B(86)) xor (A(13) and B(85)) xor (A(14) and B(84)) xor (A(15) and B(83)) xor (A(16) and B(82)) xor (A(17) and B(81)) xor (A(18) and B(80)) xor (A(19) and B(79)) xor (A(20) and B(78)) xor (A(21) and B(77)) xor (A(23) and B(76)) xor (A(23) and B(75)) xor (A(24) and B(74)) xor (A(25) and B(73)) xor (A(26) and B(72)) xor (A(27) and B(71)) xor (A(28) and B(70)) xor (A(29) and B(69)) xor (A(30) and B(68)) xor (A(31) and B(67)) xor (A(32) and B(66)) xor (A(33) and B(65)) xor (A(34) and B(64)) xor (A(35) and B(63)) xor (A(36) and B(62)) xor (A(37) and B(61)) xor (A(38) and B(60)) xor (A(39) and B(59)) xor (A(40) and B(58)) xor (A(41) and B(57)) xor (A(42) and B(56)) xor (A(43) and B(55)) xor (A(44) and B(54)) xor (A(45) and B(53)) xor (A(46) and B(52)) xor (A(47) and B(51)) xor (A(48) and B(50)) xor (A(49) and B(49)) xor (A(50) and B(48)) xor (A(51) and B(47)) xor (A(52) and B(46)) xor (A(53) and B(45)) xor (A(54) and B(44)) xor (A(55) and B(43)) xor (A(56) and B(42)) xor (A(57) and B(41)) xor (A(58) and B(40)) xor (A(59) and B(39)) xor (A(60) and B(38)) xor (A(61) and B(37)) xor (A(62) and B(36)) xor (A(63) and B(35)) xor (A(64) and B(34)) xor (A(65) and B(33)) xor (A(66) and B(32)) xor (A(67) and B(31)) xor (A(68) and B(30)) xor (A(69) and B(29)) xor (A(70) and B(28)) xor (A(71) and B(27)) xor (A(72) and B(26)) xor (A(73) and B(25)) xor (A(74) and B(24)) xor (A(75) and B(23)) xor (A(76) and B(23)) xor (A(77) and B(21)) xor (A(78) and B(20)) xor (A(79) and B(19)) xor (A(80) and B(18)) xor (A(81) and B(17)) xor (A(82) and B(16)) xor (A(83) and B(15)) xor (A(84) and B(14)) xor (A(85) and B(13)) xor (A(86) and B(12)) xor (A(87) and B(11)) xor (A(88) and B(10)) xor (A(89) and B(9)) xor (A(90) and B(8)) xor (A(91) and B(7)) xor (A(92) and B(6)) xor (A(93) and B(5)) xor (A(94) and B(4)) xor (A(95) and B(3)) xor (A(96) and B(2)) xor (A(97) and B(1)) xor (A(98) and B(0)) xor (A(91) and B(127)) xor (A(92) and B(126)) xor (A(93) and B(125)) xor (A(94) and B(124)) xor (A(95) and B(123)) xor (A(96) and B(122)) xor (A(97) and B(121)) xor (A(98) and B(120)) xor (A(99) and B(119)) xor (A(100) and B(118)) xor (A(101) and B(117)) xor (A(102) and B(116)) xor (A(103) and B(115)) xor (A(104) and B(114)) xor (A(105) and B(113)) xor (A(106) and B(112)) xor (A(107) and B(111)) xor (A(108) and B(110)) xor (A(109) and B(109)) xor (A(110) and B(108)) xor (A(111) and B(107)) xor (A(112) and B(106)) xor (A(113) and B(105)) xor (A(114) and B(104)) xor (A(115) and B(103)) xor (A(116) and B(102)) xor (A(117) and B(101)) xor (A(118) and B(100)) xor (A(119) and B(99)) xor (A(120) and B(98)) xor (A(121) and B(97)) xor (A(122) and B(96)) xor (A(123) and B(95)) xor (A(124) and B(94)) xor (A(125) and B(93)) xor (A(126) and B(92)) xor (A(96) and B(127)) xor (A(97) and B(126)) xor (A(98) and B(125)) xor (A(99) and B(124)) xor (A(100) and B(123)) xor (A(101) and B(122)) xor (A(102) and B(121)) xor (A(103) and B(120)) xor (A(104) and B(119)) xor (A(105) and B(118)) xor (A(106) and B(117)) xor (A(107) and B(116)) xor (A(108) and B(115)) xor (A(109) and B(114)) xor (A(110) and B(113)) xor (A(111) and B(112)) xor (A(112) and B(111)) xor (A(113) and B(110)) xor (A(114) and B(109)) xor (A(115) and B(108)) xor (A(116) and B(107)) xor (A(117) and B(106)) xor (A(118) and B(105)) xor (A(119) and B(104)) xor (A(120) and B(103)) xor (A(121) and B(102)) xor (A(122) and B(101)) xor (A(123) and B(100)) xor (A(124) and B(99)) xor (A(125) and B(98)) xor (A(126) and B(97)) xor (A(97) and B(127)) xor (A(98) and B(126)) xor (A(99) and B(125)) xor (A(100) and B(124)) xor (A(101) and B(123)) xor (A(102) and B(122)) xor (A(103) and B(121)) xor (A(104) and B(120)) xor (A(105) and B(119)) xor (A(106) and B(118)) xor (A(107) and B(117)) xor (A(108) and B(116)) xor (A(109) and B(115)) xor (A(110) and B(114)) xor (A(111) and B(113)) xor (A(112) and B(112)) xor (A(113) and B(111)) xor (A(114) and B(110)) xor (A(115) and B(109)) xor (A(116) and B(108)) xor (A(117) and B(107)) xor (A(118) and B(106)) xor (A(119) and B(105)) xor (A(120) and B(104)) xor (A(121) and B(103)) xor (A(122) and B(102)) xor (A(123) and B(101)) xor (A(124) and B(100)) xor (A(125) and B(99)) xor (A(126) and B(98)) xor (A(98) and B(127)) xor (A(99) and B(126)) xor (A(100) and B(125)) xor (A(101) and B(124)) xor (A(102) and B(123)) xor (A(103) and B(122)) xor (A(104) and B(121)) xor (A(105) and B(120)) xor (A(106) and B(119)) xor (A(107) and B(118)) xor (A(108) and B(117)) xor (A(109) and B(116)) xor (A(110) and B(115)) xor (A(111) and B(114)) xor (A(112) and B(113)) xor (A(113) and B(112)) xor (A(114) and B(111)) xor (A(115) and B(110)) xor (A(116) and B(109)) xor (A(117) and B(108)) xor (A(118) and B(107)) xor (A(119) and B(106)) xor (A(120) and B(105)) xor (A(121) and B(104)) xor (A(122) and B(103)) xor (A(123) and B(102)) xor (A(124) and B(101)) xor (A(125) and B(100)) xor (A(126) and B(100));
    C(99)  <= (A(0) and B(99)) xor (A(1) and B(98)) xor (A(2) and B(97)) xor (A(3) and B(96)) xor (A(4) and B(95)) xor (A(5) and B(94)) xor (A(6) and B(93)) xor (A(7) and B(92)) xor (A(8) and B(91)) xor (A(9) and B(90)) xor (A(10) and B(89)) xor (A(11) and B(88)) xor (A(12) and B(87)) xor (A(13) and B(86)) xor (A(14) and B(85)) xor (A(15) and B(84)) xor (A(16) and B(83)) xor (A(17) and B(82)) xor (A(18) and B(81)) xor (A(19) and B(80)) xor (A(20) and B(79)) xor (A(21) and B(78)) xor (A(23) and B(77)) xor (A(23) and B(76)) xor (A(24) and B(75)) xor (A(25) and B(74)) xor (A(26) and B(73)) xor (A(27) and B(72)) xor (A(28) and B(71)) xor (A(29) and B(70)) xor (A(30) and B(69)) xor (A(31) and B(68)) xor (A(32) and B(67)) xor (A(33) and B(66)) xor (A(34) and B(65)) xor (A(35) and B(64)) xor (A(36) and B(63)) xor (A(37) and B(62)) xor (A(38) and B(61)) xor (A(39) and B(60)) xor (A(40) and B(59)) xor (A(41) and B(58)) xor (A(42) and B(57)) xor (A(43) and B(56)) xor (A(44) and B(55)) xor (A(45) and B(54)) xor (A(46) and B(53)) xor (A(47) and B(52)) xor (A(48) and B(51)) xor (A(49) and B(50)) xor (A(50) and B(49)) xor (A(51) and B(48)) xor (A(52) and B(47)) xor (A(53) and B(46)) xor (A(54) and B(45)) xor (A(55) and B(44)) xor (A(56) and B(43)) xor (A(57) and B(42)) xor (A(58) and B(41)) xor (A(59) and B(40)) xor (A(60) and B(39)) xor (A(61) and B(38)) xor (A(62) and B(37)) xor (A(63) and B(36)) xor (A(64) and B(35)) xor (A(65) and B(34)) xor (A(66) and B(33)) xor (A(67) and B(32)) xor (A(68) and B(31)) xor (A(69) and B(30)) xor (A(70) and B(29)) xor (A(71) and B(28)) xor (A(72) and B(27)) xor (A(73) and B(26)) xor (A(74) and B(25)) xor (A(75) and B(24)) xor (A(76) and B(23)) xor (A(77) and B(23)) xor (A(78) and B(21)) xor (A(79) and B(20)) xor (A(80) and B(19)) xor (A(81) and B(18)) xor (A(82) and B(17)) xor (A(83) and B(16)) xor (A(84) and B(15)) xor (A(85) and B(14)) xor (A(86) and B(13)) xor (A(87) and B(12)) xor (A(88) and B(11)) xor (A(89) and B(10)) xor (A(90) and B(9)) xor (A(91) and B(8)) xor (A(92) and B(7)) xor (A(93) and B(6)) xor (A(94) and B(5)) xor (A(95) and B(4)) xor (A(96) and B(3)) xor (A(97) and B(2)) xor (A(98) and B(1)) xor (A(99) and B(0)) xor (A(92) and B(127)) xor (A(93) and B(126)) xor (A(94) and B(125)) xor (A(95) and B(124)) xor (A(96) and B(123)) xor (A(97) and B(122)) xor (A(98) and B(121)) xor (A(99) and B(120)) xor (A(100) and B(119)) xor (A(101) and B(118)) xor (A(102) and B(117)) xor (A(103) and B(116)) xor (A(104) and B(115)) xor (A(105) and B(114)) xor (A(106) and B(113)) xor (A(107) and B(112)) xor (A(108) and B(111)) xor (A(109) and B(110)) xor (A(110) and B(109)) xor (A(111) and B(108)) xor (A(112) and B(107)) xor (A(113) and B(106)) xor (A(114) and B(105)) xor (A(115) and B(104)) xor (A(116) and B(103)) xor (A(117) and B(102)) xor (A(118) and B(101)) xor (A(119) and B(100)) xor (A(120) and B(99)) xor (A(121) and B(98)) xor (A(122) and B(97)) xor (A(123) and B(96)) xor (A(124) and B(95)) xor (A(125) and B(94)) xor (A(126) and B(93)) xor (A(97) and B(127)) xor (A(98) and B(126)) xor (A(99) and B(125)) xor (A(100) and B(124)) xor (A(101) and B(123)) xor (A(102) and B(122)) xor (A(103) and B(121)) xor (A(104) and B(120)) xor (A(105) and B(119)) xor (A(106) and B(118)) xor (A(107) and B(117)) xor (A(108) and B(116)) xor (A(109) and B(115)) xor (A(110) and B(114)) xor (A(111) and B(113)) xor (A(112) and B(112)) xor (A(113) and B(111)) xor (A(114) and B(110)) xor (A(115) and B(109)) xor (A(116) and B(108)) xor (A(117) and B(107)) xor (A(118) and B(106)) xor (A(119) and B(105)) xor (A(120) and B(104)) xor (A(121) and B(103)) xor (A(122) and B(102)) xor (A(123) and B(101)) xor (A(124) and B(100)) xor (A(125) and B(99)) xor (A(126) and B(98)) xor (A(98) and B(127)) xor (A(99) and B(126)) xor (A(100) and B(125)) xor (A(101) and B(124)) xor (A(102) and B(123)) xor (A(103) and B(122)) xor (A(104) and B(121)) xor (A(105) and B(120)) xor (A(106) and B(119)) xor (A(107) and B(118)) xor (A(108) and B(117)) xor (A(109) and B(116)) xor (A(110) and B(115)) xor (A(111) and B(114)) xor (A(112) and B(113)) xor (A(113) and B(112)) xor (A(114) and B(111)) xor (A(115) and B(110)) xor (A(116) and B(109)) xor (A(117) and B(108)) xor (A(118) and B(107)) xor (A(119) and B(106)) xor (A(120) and B(105)) xor (A(121) and B(104)) xor (A(122) and B(103)) xor (A(123) and B(102)) xor (A(124) and B(101)) xor (A(125) and B(100)) xor (A(126) and B(99)) xor (A(99) and B(127)) xor (A(100) and B(126)) xor (A(101) and B(125)) xor (A(102) and B(124)) xor (A(103) and B(123)) xor (A(104) and B(122)) xor (A(105) and B(121)) xor (A(106) and B(120)) xor (A(107) and B(119)) xor (A(108) and B(118)) xor (A(109) and B(117)) xor (A(110) and B(116)) xor (A(111) and B(115)) xor (A(112) and B(114)) xor (A(113) and B(113)) xor (A(114) and B(112)) xor (A(115) and B(111)) xor (A(116) and B(110)) xor (A(117) and B(109)) xor (A(118) and B(108)) xor (A(119) and B(107)) xor (A(120) and B(106)) xor (A(121) and B(105)) xor (A(122) and B(104)) xor (A(123) and B(103)) xor (A(124) and B(102)) xor (A(125) and B(101)) xor (A(126) and B(101));
    C(100) <= (A(0) and B(100)) xor (A(1) and B(99)) xor (A(2) and B(98)) xor (A(3) and B(97)) xor (A(4) and B(96)) xor (A(5) and B(95)) xor (A(6) and B(94)) xor (A(7) and B(93)) xor (A(8) and B(92)) xor (A(9) and B(91)) xor (A(10) and B(90)) xor (A(11) and B(89)) xor (A(12) and B(88)) xor (A(13) and B(87)) xor (A(14) and B(86)) xor (A(15) and B(85)) xor (A(16) and B(84)) xor (A(17) and B(83)) xor (A(18) and B(82)) xor (A(19) and B(81)) xor (A(20) and B(80)) xor (A(21) and B(79)) xor (A(23) and B(78)) xor (A(23) and B(77)) xor (A(24) and B(76)) xor (A(25) and B(75)) xor (A(26) and B(74)) xor (A(27) and B(73)) xor (A(28) and B(72)) xor (A(29) and B(71)) xor (A(30) and B(70)) xor (A(31) and B(69)) xor (A(32) and B(68)) xor (A(33) and B(67)) xor (A(34) and B(66)) xor (A(35) and B(65)) xor (A(36) and B(64)) xor (A(37) and B(63)) xor (A(38) and B(62)) xor (A(39) and B(61)) xor (A(40) and B(60)) xor (A(41) and B(59)) xor (A(42) and B(58)) xor (A(43) and B(57)) xor (A(44) and B(56)) xor (A(45) and B(55)) xor (A(46) and B(54)) xor (A(47) and B(53)) xor (A(48) and B(52)) xor (A(49) and B(51)) xor (A(50) and B(50)) xor (A(51) and B(49)) xor (A(52) and B(48)) xor (A(53) and B(47)) xor (A(54) and B(46)) xor (A(55) and B(45)) xor (A(56) and B(44)) xor (A(57) and B(43)) xor (A(58) and B(42)) xor (A(59) and B(41)) xor (A(60) and B(40)) xor (A(61) and B(39)) xor (A(62) and B(38)) xor (A(63) and B(37)) xor (A(64) and B(36)) xor (A(65) and B(35)) xor (A(66) and B(34)) xor (A(67) and B(33)) xor (A(68) and B(32)) xor (A(69) and B(31)) xor (A(70) and B(30)) xor (A(71) and B(29)) xor (A(72) and B(28)) xor (A(73) and B(27)) xor (A(74) and B(26)) xor (A(75) and B(25)) xor (A(76) and B(24)) xor (A(77) and B(23)) xor (A(78) and B(23)) xor (A(79) and B(21)) xor (A(80) and B(20)) xor (A(81) and B(19)) xor (A(82) and B(18)) xor (A(83) and B(17)) xor (A(84) and B(16)) xor (A(85) and B(15)) xor (A(86) and B(14)) xor (A(87) and B(13)) xor (A(88) and B(12)) xor (A(89) and B(11)) xor (A(90) and B(10)) xor (A(91) and B(9)) xor (A(92) and B(8)) xor (A(93) and B(7)) xor (A(94) and B(6)) xor (A(95) and B(5)) xor (A(96) and B(4)) xor (A(97) and B(3)) xor (A(98) and B(2)) xor (A(99) and B(1)) xor (A(100) and B(0)) xor (A(93) and B(127)) xor (A(94) and B(126)) xor (A(95) and B(125)) xor (A(96) and B(124)) xor (A(97) and B(123)) xor (A(98) and B(122)) xor (A(99) and B(121)) xor (A(100) and B(120)) xor (A(101) and B(119)) xor (A(102) and B(118)) xor (A(103) and B(117)) xor (A(104) and B(116)) xor (A(105) and B(115)) xor (A(106) and B(114)) xor (A(107) and B(113)) xor (A(108) and B(112)) xor (A(109) and B(111)) xor (A(110) and B(110)) xor (A(111) and B(109)) xor (A(112) and B(108)) xor (A(113) and B(107)) xor (A(114) and B(106)) xor (A(115) and B(105)) xor (A(116) and B(104)) xor (A(117) and B(103)) xor (A(118) and B(102)) xor (A(119) and B(101)) xor (A(120) and B(100)) xor (A(121) and B(99)) xor (A(122) and B(98)) xor (A(123) and B(97)) xor (A(124) and B(96)) xor (A(125) and B(95)) xor (A(126) and B(94)) xor (A(98) and B(127)) xor (A(99) and B(126)) xor (A(100) and B(125)) xor (A(101) and B(124)) xor (A(102) and B(123)) xor (A(103) and B(122)) xor (A(104) and B(121)) xor (A(105) and B(120)) xor (A(106) and B(119)) xor (A(107) and B(118)) xor (A(108) and B(117)) xor (A(109) and B(116)) xor (A(110) and B(115)) xor (A(111) and B(114)) xor (A(112) and B(113)) xor (A(113) and B(112)) xor (A(114) and B(111)) xor (A(115) and B(110)) xor (A(116) and B(109)) xor (A(117) and B(108)) xor (A(118) and B(107)) xor (A(119) and B(106)) xor (A(120) and B(105)) xor (A(121) and B(104)) xor (A(122) and B(103)) xor (A(123) and B(102)) xor (A(124) and B(101)) xor (A(125) and B(100)) xor (A(126) and B(99)) xor (A(99) and B(127)) xor (A(100) and B(126)) xor (A(101) and B(125)) xor (A(102) and B(124)) xor (A(103) and B(123)) xor (A(104) and B(122)) xor (A(105) and B(121)) xor (A(106) and B(120)) xor (A(107) and B(119)) xor (A(108) and B(118)) xor (A(109) and B(117)) xor (A(110) and B(116)) xor (A(111) and B(115)) xor (A(112) and B(114)) xor (A(113) and B(113)) xor (A(114) and B(112)) xor (A(115) and B(111)) xor (A(116) and B(110)) xor (A(117) and B(109)) xor (A(118) and B(108)) xor (A(119) and B(107)) xor (A(120) and B(106)) xor (A(121) and B(105)) xor (A(122) and B(104)) xor (A(123) and B(103)) xor (A(124) and B(102)) xor (A(125) and B(101)) xor (A(126) and B(100)) xor (A(100) and B(127)) xor (A(101) and B(126)) xor (A(102) and B(125)) xor (A(103) and B(124)) xor (A(104) and B(123)) xor (A(105) and B(122)) xor (A(106) and B(121)) xor (A(107) and B(120)) xor (A(108) and B(119)) xor (A(109) and B(118)) xor (A(110) and B(117)) xor (A(111) and B(116)) xor (A(112) and B(115)) xor (A(113) and B(114)) xor (A(114) and B(113)) xor (A(115) and B(112)) xor (A(116) and B(111)) xor (A(117) and B(110)) xor (A(118) and B(109)) xor (A(119) and B(108)) xor (A(120) and B(107)) xor (A(121) and B(106)) xor (A(122) and B(105)) xor (A(123) and B(104)) xor (A(124) and B(103)) xor (A(125) and B(102)) xor (A(126) and B(102));
    C(101) <= (A(0) and B(101)) xor (A(1) and B(100)) xor (A(2) and B(99)) xor (A(3) and B(98)) xor (A(4) and B(97)) xor (A(5) and B(96)) xor (A(6) and B(95)) xor (A(7) and B(94)) xor (A(8) and B(93)) xor (A(9) and B(92)) xor (A(10) and B(91)) xor (A(11) and B(90)) xor (A(12) and B(89)) xor (A(13) and B(88)) xor (A(14) and B(87)) xor (A(15) and B(86)) xor (A(16) and B(85)) xor (A(17) and B(84)) xor (A(18) and B(83)) xor (A(19) and B(82)) xor (A(20) and B(81)) xor (A(21) and B(80)) xor (A(23) and B(79)) xor (A(23) and B(78)) xor (A(24) and B(77)) xor (A(25) and B(76)) xor (A(26) and B(75)) xor (A(27) and B(74)) xor (A(28) and B(73)) xor (A(29) and B(72)) xor (A(30) and B(71)) xor (A(31) and B(70)) xor (A(32) and B(69)) xor (A(33) and B(68)) xor (A(34) and B(67)) xor (A(35) and B(66)) xor (A(36) and B(65)) xor (A(37) and B(64)) xor (A(38) and B(63)) xor (A(39) and B(62)) xor (A(40) and B(61)) xor (A(41) and B(60)) xor (A(42) and B(59)) xor (A(43) and B(58)) xor (A(44) and B(57)) xor (A(45) and B(56)) xor (A(46) and B(55)) xor (A(47) and B(54)) xor (A(48) and B(53)) xor (A(49) and B(52)) xor (A(50) and B(51)) xor (A(51) and B(50)) xor (A(52) and B(49)) xor (A(53) and B(48)) xor (A(54) and B(47)) xor (A(55) and B(46)) xor (A(56) and B(45)) xor (A(57) and B(44)) xor (A(58) and B(43)) xor (A(59) and B(42)) xor (A(60) and B(41)) xor (A(61) and B(40)) xor (A(62) and B(39)) xor (A(63) and B(38)) xor (A(64) and B(37)) xor (A(65) and B(36)) xor (A(66) and B(35)) xor (A(67) and B(34)) xor (A(68) and B(33)) xor (A(69) and B(32)) xor (A(70) and B(31)) xor (A(71) and B(30)) xor (A(72) and B(29)) xor (A(73) and B(28)) xor (A(74) and B(27)) xor (A(75) and B(26)) xor (A(76) and B(25)) xor (A(77) and B(24)) xor (A(78) and B(23)) xor (A(79) and B(23)) xor (A(80) and B(21)) xor (A(81) and B(20)) xor (A(82) and B(19)) xor (A(83) and B(18)) xor (A(84) and B(17)) xor (A(85) and B(16)) xor (A(86) and B(15)) xor (A(87) and B(14)) xor (A(88) and B(13)) xor (A(89) and B(12)) xor (A(90) and B(11)) xor (A(91) and B(10)) xor (A(92) and B(9)) xor (A(93) and B(8)) xor (A(94) and B(7)) xor (A(95) and B(6)) xor (A(96) and B(5)) xor (A(97) and B(4)) xor (A(98) and B(3)) xor (A(99) and B(2)) xor (A(100) and B(1)) xor (A(101) and B(0)) xor (A(94) and B(127)) xor (A(95) and B(126)) xor (A(96) and B(125)) xor (A(97) and B(124)) xor (A(98) and B(123)) xor (A(99) and B(122)) xor (A(100) and B(121)) xor (A(101) and B(120)) xor (A(102) and B(119)) xor (A(103) and B(118)) xor (A(104) and B(117)) xor (A(105) and B(116)) xor (A(106) and B(115)) xor (A(107) and B(114)) xor (A(108) and B(113)) xor (A(109) and B(112)) xor (A(110) and B(111)) xor (A(111) and B(110)) xor (A(112) and B(109)) xor (A(113) and B(108)) xor (A(114) and B(107)) xor (A(115) and B(106)) xor (A(116) and B(105)) xor (A(117) and B(104)) xor (A(118) and B(103)) xor (A(119) and B(102)) xor (A(120) and B(101)) xor (A(121) and B(100)) xor (A(122) and B(99)) xor (A(123) and B(98)) xor (A(124) and B(97)) xor (A(125) and B(96)) xor (A(126) and B(95)) xor (A(99) and B(127)) xor (A(100) and B(126)) xor (A(101) and B(125)) xor (A(102) and B(124)) xor (A(103) and B(123)) xor (A(104) and B(122)) xor (A(105) and B(121)) xor (A(106) and B(120)) xor (A(107) and B(119)) xor (A(108) and B(118)) xor (A(109) and B(117)) xor (A(110) and B(116)) xor (A(111) and B(115)) xor (A(112) and B(114)) xor (A(113) and B(113)) xor (A(114) and B(112)) xor (A(115) and B(111)) xor (A(116) and B(110)) xor (A(117) and B(109)) xor (A(118) and B(108)) xor (A(119) and B(107)) xor (A(120) and B(106)) xor (A(121) and B(105)) xor (A(122) and B(104)) xor (A(123) and B(103)) xor (A(124) and B(102)) xor (A(125) and B(101)) xor (A(126) and B(100)) xor (A(100) and B(127)) xor (A(101) and B(126)) xor (A(102) and B(125)) xor (A(103) and B(124)) xor (A(104) and B(123)) xor (A(105) and B(122)) xor (A(106) and B(121)) xor (A(107) and B(120)) xor (A(108) and B(119)) xor (A(109) and B(118)) xor (A(110) and B(117)) xor (A(111) and B(116)) xor (A(112) and B(115)) xor (A(113) and B(114)) xor (A(114) and B(113)) xor (A(115) and B(112)) xor (A(116) and B(111)) xor (A(117) and B(110)) xor (A(118) and B(109)) xor (A(119) and B(108)) xor (A(120) and B(107)) xor (A(121) and B(106)) xor (A(122) and B(105)) xor (A(123) and B(104)) xor (A(124) and B(103)) xor (A(125) and B(102)) xor (A(126) and B(101)) xor (A(101) and B(127)) xor (A(102) and B(126)) xor (A(103) and B(125)) xor (A(104) and B(124)) xor (A(105) and B(123)) xor (A(106) and B(122)) xor (A(107) and B(121)) xor (A(108) and B(120)) xor (A(109) and B(119)) xor (A(110) and B(118)) xor (A(111) and B(117)) xor (A(112) and B(116)) xor (A(113) and B(115)) xor (A(114) and B(114)) xor (A(115) and B(113)) xor (A(116) and B(112)) xor (A(117) and B(111)) xor (A(118) and B(110)) xor (A(119) and B(109)) xor (A(120) and B(108)) xor (A(121) and B(107)) xor (A(122) and B(106)) xor (A(123) and B(105)) xor (A(124) and B(104)) xor (A(125) and B(103)) xor (A(126) and B(103));
    C(102) <= (A(0) and B(102)) xor (A(1) and B(101)) xor (A(2) and B(100)) xor (A(3) and B(99)) xor (A(4) and B(98)) xor (A(5) and B(97)) xor (A(6) and B(96)) xor (A(7) and B(95)) xor (A(8) and B(94)) xor (A(9) and B(93)) xor (A(10) and B(92)) xor (A(11) and B(91)) xor (A(12) and B(90)) xor (A(13) and B(89)) xor (A(14) and B(88)) xor (A(15) and B(87)) xor (A(16) and B(86)) xor (A(17) and B(85)) xor (A(18) and B(84)) xor (A(19) and B(83)) xor (A(20) and B(82)) xor (A(21) and B(81)) xor (A(23) and B(80)) xor (A(23) and B(79)) xor (A(24) and B(78)) xor (A(25) and B(77)) xor (A(26) and B(76)) xor (A(27) and B(75)) xor (A(28) and B(74)) xor (A(29) and B(73)) xor (A(30) and B(72)) xor (A(31) and B(71)) xor (A(32) and B(70)) xor (A(33) and B(69)) xor (A(34) and B(68)) xor (A(35) and B(67)) xor (A(36) and B(66)) xor (A(37) and B(65)) xor (A(38) and B(64)) xor (A(39) and B(63)) xor (A(40) and B(62)) xor (A(41) and B(61)) xor (A(42) and B(60)) xor (A(43) and B(59)) xor (A(44) and B(58)) xor (A(45) and B(57)) xor (A(46) and B(56)) xor (A(47) and B(55)) xor (A(48) and B(54)) xor (A(49) and B(53)) xor (A(50) and B(52)) xor (A(51) and B(51)) xor (A(52) and B(50)) xor (A(53) and B(49)) xor (A(54) and B(48)) xor (A(55) and B(47)) xor (A(56) and B(46)) xor (A(57) and B(45)) xor (A(58) and B(44)) xor (A(59) and B(43)) xor (A(60) and B(42)) xor (A(61) and B(41)) xor (A(62) and B(40)) xor (A(63) and B(39)) xor (A(64) and B(38)) xor (A(65) and B(37)) xor (A(66) and B(36)) xor (A(67) and B(35)) xor (A(68) and B(34)) xor (A(69) and B(33)) xor (A(70) and B(32)) xor (A(71) and B(31)) xor (A(72) and B(30)) xor (A(73) and B(29)) xor (A(74) and B(28)) xor (A(75) and B(27)) xor (A(76) and B(26)) xor (A(77) and B(25)) xor (A(78) and B(24)) xor (A(79) and B(23)) xor (A(80) and B(23)) xor (A(81) and B(21)) xor (A(82) and B(20)) xor (A(83) and B(19)) xor (A(84) and B(18)) xor (A(85) and B(17)) xor (A(86) and B(16)) xor (A(87) and B(15)) xor (A(88) and B(14)) xor (A(89) and B(13)) xor (A(90) and B(12)) xor (A(91) and B(11)) xor (A(92) and B(10)) xor (A(93) and B(9)) xor (A(94) and B(8)) xor (A(95) and B(7)) xor (A(96) and B(6)) xor (A(97) and B(5)) xor (A(98) and B(4)) xor (A(99) and B(3)) xor (A(100) and B(2)) xor (A(101) and B(1)) xor (A(102) and B(0)) xor (A(95) and B(127)) xor (A(96) and B(126)) xor (A(97) and B(125)) xor (A(98) and B(124)) xor (A(99) and B(123)) xor (A(100) and B(122)) xor (A(101) and B(121)) xor (A(102) and B(120)) xor (A(103) and B(119)) xor (A(104) and B(118)) xor (A(105) and B(117)) xor (A(106) and B(116)) xor (A(107) and B(115)) xor (A(108) and B(114)) xor (A(109) and B(113)) xor (A(110) and B(112)) xor (A(111) and B(111)) xor (A(112) and B(110)) xor (A(113) and B(109)) xor (A(114) and B(108)) xor (A(115) and B(107)) xor (A(116) and B(106)) xor (A(117) and B(105)) xor (A(118) and B(104)) xor (A(119) and B(103)) xor (A(120) and B(102)) xor (A(121) and B(101)) xor (A(122) and B(100)) xor (A(123) and B(99)) xor (A(124) and B(98)) xor (A(125) and B(97)) xor (A(126) and B(96)) xor (A(100) and B(127)) xor (A(101) and B(126)) xor (A(102) and B(125)) xor (A(103) and B(124)) xor (A(104) and B(123)) xor (A(105) and B(122)) xor (A(106) and B(121)) xor (A(107) and B(120)) xor (A(108) and B(119)) xor (A(109) and B(118)) xor (A(110) and B(117)) xor (A(111) and B(116)) xor (A(112) and B(115)) xor (A(113) and B(114)) xor (A(114) and B(113)) xor (A(115) and B(112)) xor (A(116) and B(111)) xor (A(117) and B(110)) xor (A(118) and B(109)) xor (A(119) and B(108)) xor (A(120) and B(107)) xor (A(121) and B(106)) xor (A(122) and B(105)) xor (A(123) and B(104)) xor (A(124) and B(103)) xor (A(125) and B(102)) xor (A(126) and B(101)) xor (A(101) and B(127)) xor (A(102) and B(126)) xor (A(103) and B(125)) xor (A(104) and B(124)) xor (A(105) and B(123)) xor (A(106) and B(122)) xor (A(107) and B(121)) xor (A(108) and B(120)) xor (A(109) and B(119)) xor (A(110) and B(118)) xor (A(111) and B(117)) xor (A(112) and B(116)) xor (A(113) and B(115)) xor (A(114) and B(114)) xor (A(115) and B(113)) xor (A(116) and B(112)) xor (A(117) and B(111)) xor (A(118) and B(110)) xor (A(119) and B(109)) xor (A(120) and B(108)) xor (A(121) and B(107)) xor (A(122) and B(106)) xor (A(123) and B(105)) xor (A(124) and B(104)) xor (A(125) and B(103)) xor (A(126) and B(102)) xor (A(102) and B(127)) xor (A(103) and B(126)) xor (A(104) and B(125)) xor (A(105) and B(124)) xor (A(106) and B(123)) xor (A(107) and B(122)) xor (A(108) and B(121)) xor (A(109) and B(120)) xor (A(110) and B(119)) xor (A(111) and B(118)) xor (A(112) and B(117)) xor (A(113) and B(116)) xor (A(114) and B(115)) xor (A(115) and B(114)) xor (A(116) and B(113)) xor (A(117) and B(112)) xor (A(118) and B(111)) xor (A(119) and B(110)) xor (A(120) and B(109)) xor (A(121) and B(108)) xor (A(122) and B(107)) xor (A(123) and B(106)) xor (A(124) and B(105)) xor (A(125) and B(104)) xor (A(126) and B(104));
    C(103) <= (A(0) and B(103)) xor (A(1) and B(102)) xor (A(2) and B(101)) xor (A(3) and B(100)) xor (A(4) and B(99)) xor (A(5) and B(98)) xor (A(6) and B(97)) xor (A(7) and B(96)) xor (A(8) and B(95)) xor (A(9) and B(94)) xor (A(10) and B(93)) xor (A(11) and B(92)) xor (A(12) and B(91)) xor (A(13) and B(90)) xor (A(14) and B(89)) xor (A(15) and B(88)) xor (A(16) and B(87)) xor (A(17) and B(86)) xor (A(18) and B(85)) xor (A(19) and B(84)) xor (A(20) and B(83)) xor (A(21) and B(82)) xor (A(23) and B(81)) xor (A(23) and B(80)) xor (A(24) and B(79)) xor (A(25) and B(78)) xor (A(26) and B(77)) xor (A(27) and B(76)) xor (A(28) and B(75)) xor (A(29) and B(74)) xor (A(30) and B(73)) xor (A(31) and B(72)) xor (A(32) and B(71)) xor (A(33) and B(70)) xor (A(34) and B(69)) xor (A(35) and B(68)) xor (A(36) and B(67)) xor (A(37) and B(66)) xor (A(38) and B(65)) xor (A(39) and B(64)) xor (A(40) and B(63)) xor (A(41) and B(62)) xor (A(42) and B(61)) xor (A(43) and B(60)) xor (A(44) and B(59)) xor (A(45) and B(58)) xor (A(46) and B(57)) xor (A(47) and B(56)) xor (A(48) and B(55)) xor (A(49) and B(54)) xor (A(50) and B(53)) xor (A(51) and B(52)) xor (A(52) and B(51)) xor (A(53) and B(50)) xor (A(54) and B(49)) xor (A(55) and B(48)) xor (A(56) and B(47)) xor (A(57) and B(46)) xor (A(58) and B(45)) xor (A(59) and B(44)) xor (A(60) and B(43)) xor (A(61) and B(42)) xor (A(62) and B(41)) xor (A(63) and B(40)) xor (A(64) and B(39)) xor (A(65) and B(38)) xor (A(66) and B(37)) xor (A(67) and B(36)) xor (A(68) and B(35)) xor (A(69) and B(34)) xor (A(70) and B(33)) xor (A(71) and B(32)) xor (A(72) and B(31)) xor (A(73) and B(30)) xor (A(74) and B(29)) xor (A(75) and B(28)) xor (A(76) and B(27)) xor (A(77) and B(26)) xor (A(78) and B(25)) xor (A(79) and B(24)) xor (A(80) and B(23)) xor (A(81) and B(23)) xor (A(82) and B(21)) xor (A(83) and B(20)) xor (A(84) and B(19)) xor (A(85) and B(18)) xor (A(86) and B(17)) xor (A(87) and B(16)) xor (A(88) and B(15)) xor (A(89) and B(14)) xor (A(90) and B(13)) xor (A(91) and B(12)) xor (A(92) and B(11)) xor (A(93) and B(10)) xor (A(94) and B(9)) xor (A(95) and B(8)) xor (A(96) and B(7)) xor (A(97) and B(6)) xor (A(98) and B(5)) xor (A(99) and B(4)) xor (A(100) and B(3)) xor (A(101) and B(2)) xor (A(102) and B(1)) xor (A(103) and B(0)) xor (A(96) and B(127)) xor (A(97) and B(126)) xor (A(98) and B(125)) xor (A(99) and B(124)) xor (A(100) and B(123)) xor (A(101) and B(122)) xor (A(102) and B(121)) xor (A(103) and B(120)) xor (A(104) and B(119)) xor (A(105) and B(118)) xor (A(106) and B(117)) xor (A(107) and B(116)) xor (A(108) and B(115)) xor (A(109) and B(114)) xor (A(110) and B(113)) xor (A(111) and B(112)) xor (A(112) and B(111)) xor (A(113) and B(110)) xor (A(114) and B(109)) xor (A(115) and B(108)) xor (A(116) and B(107)) xor (A(117) and B(106)) xor (A(118) and B(105)) xor (A(119) and B(104)) xor (A(120) and B(103)) xor (A(121) and B(102)) xor (A(122) and B(101)) xor (A(123) and B(100)) xor (A(124) and B(99)) xor (A(125) and B(98)) xor (A(126) and B(97)) xor (A(101) and B(127)) xor (A(102) and B(126)) xor (A(103) and B(125)) xor (A(104) and B(124)) xor (A(105) and B(123)) xor (A(106) and B(122)) xor (A(107) and B(121)) xor (A(108) and B(120)) xor (A(109) and B(119)) xor (A(110) and B(118)) xor (A(111) and B(117)) xor (A(112) and B(116)) xor (A(113) and B(115)) xor (A(114) and B(114)) xor (A(115) and B(113)) xor (A(116) and B(112)) xor (A(117) and B(111)) xor (A(118) and B(110)) xor (A(119) and B(109)) xor (A(120) and B(108)) xor (A(121) and B(107)) xor (A(122) and B(106)) xor (A(123) and B(105)) xor (A(124) and B(104)) xor (A(125) and B(103)) xor (A(126) and B(102)) xor (A(102) and B(127)) xor (A(103) and B(126)) xor (A(104) and B(125)) xor (A(105) and B(124)) xor (A(106) and B(123)) xor (A(107) and B(122)) xor (A(108) and B(121)) xor (A(109) and B(120)) xor (A(110) and B(119)) xor (A(111) and B(118)) xor (A(112) and B(117)) xor (A(113) and B(116)) xor (A(114) and B(115)) xor (A(115) and B(114)) xor (A(116) and B(113)) xor (A(117) and B(112)) xor (A(118) and B(111)) xor (A(119) and B(110)) xor (A(120) and B(109)) xor (A(121) and B(108)) xor (A(122) and B(107)) xor (A(123) and B(106)) xor (A(124) and B(105)) xor (A(125) and B(104)) xor (A(126) and B(103)) xor (A(103) and B(127)) xor (A(104) and B(126)) xor (A(105) and B(125)) xor (A(106) and B(124)) xor (A(107) and B(123)) xor (A(108) and B(122)) xor (A(109) and B(121)) xor (A(110) and B(120)) xor (A(111) and B(119)) xor (A(112) and B(118)) xor (A(113) and B(117)) xor (A(114) and B(116)) xor (A(115) and B(115)) xor (A(116) and B(114)) xor (A(117) and B(113)) xor (A(118) and B(112)) xor (A(119) and B(111)) xor (A(120) and B(110)) xor (A(121) and B(109)) xor (A(122) and B(108)) xor (A(123) and B(107)) xor (A(124) and B(106)) xor (A(125) and B(105)) xor (A(126) and B(105));
    C(104) <= (A(0) and B(104)) xor (A(1) and B(103)) xor (A(2) and B(102)) xor (A(3) and B(101)) xor (A(4) and B(100)) xor (A(5) and B(99)) xor (A(6) and B(98)) xor (A(7) and B(97)) xor (A(8) and B(96)) xor (A(9) and B(95)) xor (A(10) and B(94)) xor (A(11) and B(93)) xor (A(12) and B(92)) xor (A(13) and B(91)) xor (A(14) and B(90)) xor (A(15) and B(89)) xor (A(16) and B(88)) xor (A(17) and B(87)) xor (A(18) and B(86)) xor (A(19) and B(85)) xor (A(20) and B(84)) xor (A(21) and B(83)) xor (A(23) and B(82)) xor (A(23) and B(81)) xor (A(24) and B(80)) xor (A(25) and B(79)) xor (A(26) and B(78)) xor (A(27) and B(77)) xor (A(28) and B(76)) xor (A(29) and B(75)) xor (A(30) and B(74)) xor (A(31) and B(73)) xor (A(32) and B(72)) xor (A(33) and B(71)) xor (A(34) and B(70)) xor (A(35) and B(69)) xor (A(36) and B(68)) xor (A(37) and B(67)) xor (A(38) and B(66)) xor (A(39) and B(65)) xor (A(40) and B(64)) xor (A(41) and B(63)) xor (A(42) and B(62)) xor (A(43) and B(61)) xor (A(44) and B(60)) xor (A(45) and B(59)) xor (A(46) and B(58)) xor (A(47) and B(57)) xor (A(48) and B(56)) xor (A(49) and B(55)) xor (A(50) and B(54)) xor (A(51) and B(53)) xor (A(52) and B(52)) xor (A(53) and B(51)) xor (A(54) and B(50)) xor (A(55) and B(49)) xor (A(56) and B(48)) xor (A(57) and B(47)) xor (A(58) and B(46)) xor (A(59) and B(45)) xor (A(60) and B(44)) xor (A(61) and B(43)) xor (A(62) and B(42)) xor (A(63) and B(41)) xor (A(64) and B(40)) xor (A(65) and B(39)) xor (A(66) and B(38)) xor (A(67) and B(37)) xor (A(68) and B(36)) xor (A(69) and B(35)) xor (A(70) and B(34)) xor (A(71) and B(33)) xor (A(72) and B(32)) xor (A(73) and B(31)) xor (A(74) and B(30)) xor (A(75) and B(29)) xor (A(76) and B(28)) xor (A(77) and B(27)) xor (A(78) and B(26)) xor (A(79) and B(25)) xor (A(80) and B(24)) xor (A(81) and B(23)) xor (A(82) and B(23)) xor (A(83) and B(21)) xor (A(84) and B(20)) xor (A(85) and B(19)) xor (A(86) and B(18)) xor (A(87) and B(17)) xor (A(88) and B(16)) xor (A(89) and B(15)) xor (A(90) and B(14)) xor (A(91) and B(13)) xor (A(92) and B(12)) xor (A(93) and B(11)) xor (A(94) and B(10)) xor (A(95) and B(9)) xor (A(96) and B(8)) xor (A(97) and B(7)) xor (A(98) and B(6)) xor (A(99) and B(5)) xor (A(100) and B(4)) xor (A(101) and B(3)) xor (A(102) and B(2)) xor (A(103) and B(1)) xor (A(104) and B(0)) xor (A(97) and B(127)) xor (A(98) and B(126)) xor (A(99) and B(125)) xor (A(100) and B(124)) xor (A(101) and B(123)) xor (A(102) and B(122)) xor (A(103) and B(121)) xor (A(104) and B(120)) xor (A(105) and B(119)) xor (A(106) and B(118)) xor (A(107) and B(117)) xor (A(108) and B(116)) xor (A(109) and B(115)) xor (A(110) and B(114)) xor (A(111) and B(113)) xor (A(112) and B(112)) xor (A(113) and B(111)) xor (A(114) and B(110)) xor (A(115) and B(109)) xor (A(116) and B(108)) xor (A(117) and B(107)) xor (A(118) and B(106)) xor (A(119) and B(105)) xor (A(120) and B(104)) xor (A(121) and B(103)) xor (A(122) and B(102)) xor (A(123) and B(101)) xor (A(124) and B(100)) xor (A(125) and B(99)) xor (A(126) and B(98)) xor (A(102) and B(127)) xor (A(103) and B(126)) xor (A(104) and B(125)) xor (A(105) and B(124)) xor (A(106) and B(123)) xor (A(107) and B(122)) xor (A(108) and B(121)) xor (A(109) and B(120)) xor (A(110) and B(119)) xor (A(111) and B(118)) xor (A(112) and B(117)) xor (A(113) and B(116)) xor (A(114) and B(115)) xor (A(115) and B(114)) xor (A(116) and B(113)) xor (A(117) and B(112)) xor (A(118) and B(111)) xor (A(119) and B(110)) xor (A(120) and B(109)) xor (A(121) and B(108)) xor (A(122) and B(107)) xor (A(123) and B(106)) xor (A(124) and B(105)) xor (A(125) and B(104)) xor (A(126) and B(103)) xor (A(103) and B(127)) xor (A(104) and B(126)) xor (A(105) and B(125)) xor (A(106) and B(124)) xor (A(107) and B(123)) xor (A(108) and B(122)) xor (A(109) and B(121)) xor (A(110) and B(120)) xor (A(111) and B(119)) xor (A(112) and B(118)) xor (A(113) and B(117)) xor (A(114) and B(116)) xor (A(115) and B(115)) xor (A(116) and B(114)) xor (A(117) and B(113)) xor (A(118) and B(112)) xor (A(119) and B(111)) xor (A(120) and B(110)) xor (A(121) and B(109)) xor (A(122) and B(108)) xor (A(123) and B(107)) xor (A(124) and B(106)) xor (A(125) and B(105)) xor (A(126) and B(104)) xor (A(104) and B(127)) xor (A(105) and B(126)) xor (A(106) and B(125)) xor (A(107) and B(124)) xor (A(108) and B(123)) xor (A(109) and B(122)) xor (A(110) and B(121)) xor (A(111) and B(120)) xor (A(112) and B(119)) xor (A(113) and B(118)) xor (A(114) and B(117)) xor (A(115) and B(116)) xor (A(116) and B(115)) xor (A(117) and B(114)) xor (A(118) and B(113)) xor (A(119) and B(112)) xor (A(120) and B(111)) xor (A(121) and B(110)) xor (A(122) and B(109)) xor (A(123) and B(108)) xor (A(124) and B(107)) xor (A(125) and B(106)) xor (A(126) and B(106));
    C(105) <= (A(0) and B(105)) xor (A(1) and B(104)) xor (A(2) and B(103)) xor (A(3) and B(102)) xor (A(4) and B(101)) xor (A(5) and B(100)) xor (A(6) and B(99)) xor (A(7) and B(98)) xor (A(8) and B(97)) xor (A(9) and B(96)) xor (A(10) and B(95)) xor (A(11) and B(94)) xor (A(12) and B(93)) xor (A(13) and B(92)) xor (A(14) and B(91)) xor (A(15) and B(90)) xor (A(16) and B(89)) xor (A(17) and B(88)) xor (A(18) and B(87)) xor (A(19) and B(86)) xor (A(20) and B(85)) xor (A(21) and B(84)) xor (A(23) and B(83)) xor (A(23) and B(82)) xor (A(24) and B(81)) xor (A(25) and B(80)) xor (A(26) and B(79)) xor (A(27) and B(78)) xor (A(28) and B(77)) xor (A(29) and B(76)) xor (A(30) and B(75)) xor (A(31) and B(74)) xor (A(32) and B(73)) xor (A(33) and B(72)) xor (A(34) and B(71)) xor (A(35) and B(70)) xor (A(36) and B(69)) xor (A(37) and B(68)) xor (A(38) and B(67)) xor (A(39) and B(66)) xor (A(40) and B(65)) xor (A(41) and B(64)) xor (A(42) and B(63)) xor (A(43) and B(62)) xor (A(44) and B(61)) xor (A(45) and B(60)) xor (A(46) and B(59)) xor (A(47) and B(58)) xor (A(48) and B(57)) xor (A(49) and B(56)) xor (A(50) and B(55)) xor (A(51) and B(54)) xor (A(52) and B(53)) xor (A(53) and B(52)) xor (A(54) and B(51)) xor (A(55) and B(50)) xor (A(56) and B(49)) xor (A(57) and B(48)) xor (A(58) and B(47)) xor (A(59) and B(46)) xor (A(60) and B(45)) xor (A(61) and B(44)) xor (A(62) and B(43)) xor (A(63) and B(42)) xor (A(64) and B(41)) xor (A(65) and B(40)) xor (A(66) and B(39)) xor (A(67) and B(38)) xor (A(68) and B(37)) xor (A(69) and B(36)) xor (A(70) and B(35)) xor (A(71) and B(34)) xor (A(72) and B(33)) xor (A(73) and B(32)) xor (A(74) and B(31)) xor (A(75) and B(30)) xor (A(76) and B(29)) xor (A(77) and B(28)) xor (A(78) and B(27)) xor (A(79) and B(26)) xor (A(80) and B(25)) xor (A(81) and B(24)) xor (A(82) and B(23)) xor (A(83) and B(23)) xor (A(84) and B(21)) xor (A(85) and B(20)) xor (A(86) and B(19)) xor (A(87) and B(18)) xor (A(88) and B(17)) xor (A(89) and B(16)) xor (A(90) and B(15)) xor (A(91) and B(14)) xor (A(92) and B(13)) xor (A(93) and B(12)) xor (A(94) and B(11)) xor (A(95) and B(10)) xor (A(96) and B(9)) xor (A(97) and B(8)) xor (A(98) and B(7)) xor (A(99) and B(6)) xor (A(100) and B(5)) xor (A(101) and B(4)) xor (A(102) and B(3)) xor (A(103) and B(2)) xor (A(104) and B(1)) xor (A(105) and B(0)) xor (A(98) and B(127)) xor (A(99) and B(126)) xor (A(100) and B(125)) xor (A(101) and B(124)) xor (A(102) and B(123)) xor (A(103) and B(122)) xor (A(104) and B(121)) xor (A(105) and B(120)) xor (A(106) and B(119)) xor (A(107) and B(118)) xor (A(108) and B(117)) xor (A(109) and B(116)) xor (A(110) and B(115)) xor (A(111) and B(114)) xor (A(112) and B(113)) xor (A(113) and B(112)) xor (A(114) and B(111)) xor (A(115) and B(110)) xor (A(116) and B(109)) xor (A(117) and B(108)) xor (A(118) and B(107)) xor (A(119) and B(106)) xor (A(120) and B(105)) xor (A(121) and B(104)) xor (A(122) and B(103)) xor (A(123) and B(102)) xor (A(124) and B(101)) xor (A(125) and B(100)) xor (A(126) and B(99)) xor (A(103) and B(127)) xor (A(104) and B(126)) xor (A(105) and B(125)) xor (A(106) and B(124)) xor (A(107) and B(123)) xor (A(108) and B(122)) xor (A(109) and B(121)) xor (A(110) and B(120)) xor (A(111) and B(119)) xor (A(112) and B(118)) xor (A(113) and B(117)) xor (A(114) and B(116)) xor (A(115) and B(115)) xor (A(116) and B(114)) xor (A(117) and B(113)) xor (A(118) and B(112)) xor (A(119) and B(111)) xor (A(120) and B(110)) xor (A(121) and B(109)) xor (A(122) and B(108)) xor (A(123) and B(107)) xor (A(124) and B(106)) xor (A(125) and B(105)) xor (A(126) and B(104)) xor (A(104) and B(127)) xor (A(105) and B(126)) xor (A(106) and B(125)) xor (A(107) and B(124)) xor (A(108) and B(123)) xor (A(109) and B(122)) xor (A(110) and B(121)) xor (A(111) and B(120)) xor (A(112) and B(119)) xor (A(113) and B(118)) xor (A(114) and B(117)) xor (A(115) and B(116)) xor (A(116) and B(115)) xor (A(117) and B(114)) xor (A(118) and B(113)) xor (A(119) and B(112)) xor (A(120) and B(111)) xor (A(121) and B(110)) xor (A(122) and B(109)) xor (A(123) and B(108)) xor (A(124) and B(107)) xor (A(125) and B(106)) xor (A(126) and B(105)) xor (A(105) and B(127)) xor (A(106) and B(126)) xor (A(107) and B(125)) xor (A(108) and B(124)) xor (A(109) and B(123)) xor (A(110) and B(122)) xor (A(111) and B(121)) xor (A(112) and B(120)) xor (A(113) and B(119)) xor (A(114) and B(118)) xor (A(115) and B(117)) xor (A(116) and B(116)) xor (A(117) and B(115)) xor (A(118) and B(114)) xor (A(119) and B(113)) xor (A(120) and B(112)) xor (A(121) and B(111)) xor (A(122) and B(110)) xor (A(123) and B(109)) xor (A(124) and B(108)) xor (A(125) and B(107)) xor (A(126) and B(107));
    C(106) <= (A(0) and B(106)) xor (A(1) and B(105)) xor (A(2) and B(104)) xor (A(3) and B(103)) xor (A(4) and B(102)) xor (A(5) and B(101)) xor (A(6) and B(100)) xor (A(7) and B(99)) xor (A(8) and B(98)) xor (A(9) and B(97)) xor (A(10) and B(96)) xor (A(11) and B(95)) xor (A(12) and B(94)) xor (A(13) and B(93)) xor (A(14) and B(92)) xor (A(15) and B(91)) xor (A(16) and B(90)) xor (A(17) and B(89)) xor (A(18) and B(88)) xor (A(19) and B(87)) xor (A(20) and B(86)) xor (A(21) and B(85)) xor (A(23) and B(84)) xor (A(23) and B(83)) xor (A(24) and B(82)) xor (A(25) and B(81)) xor (A(26) and B(80)) xor (A(27) and B(79)) xor (A(28) and B(78)) xor (A(29) and B(77)) xor (A(30) and B(76)) xor (A(31) and B(75)) xor (A(32) and B(74)) xor (A(33) and B(73)) xor (A(34) and B(72)) xor (A(35) and B(71)) xor (A(36) and B(70)) xor (A(37) and B(69)) xor (A(38) and B(68)) xor (A(39) and B(67)) xor (A(40) and B(66)) xor (A(41) and B(65)) xor (A(42) and B(64)) xor (A(43) and B(63)) xor (A(44) and B(62)) xor (A(45) and B(61)) xor (A(46) and B(60)) xor (A(47) and B(59)) xor (A(48) and B(58)) xor (A(49) and B(57)) xor (A(50) and B(56)) xor (A(51) and B(55)) xor (A(52) and B(54)) xor (A(53) and B(53)) xor (A(54) and B(52)) xor (A(55) and B(51)) xor (A(56) and B(50)) xor (A(57) and B(49)) xor (A(58) and B(48)) xor (A(59) and B(47)) xor (A(60) and B(46)) xor (A(61) and B(45)) xor (A(62) and B(44)) xor (A(63) and B(43)) xor (A(64) and B(42)) xor (A(65) and B(41)) xor (A(66) and B(40)) xor (A(67) and B(39)) xor (A(68) and B(38)) xor (A(69) and B(37)) xor (A(70) and B(36)) xor (A(71) and B(35)) xor (A(72) and B(34)) xor (A(73) and B(33)) xor (A(74) and B(32)) xor (A(75) and B(31)) xor (A(76) and B(30)) xor (A(77) and B(29)) xor (A(78) and B(28)) xor (A(79) and B(27)) xor (A(80) and B(26)) xor (A(81) and B(25)) xor (A(82) and B(24)) xor (A(83) and B(23)) xor (A(84) and B(23)) xor (A(85) and B(21)) xor (A(86) and B(20)) xor (A(87) and B(19)) xor (A(88) and B(18)) xor (A(89) and B(17)) xor (A(90) and B(16)) xor (A(91) and B(15)) xor (A(92) and B(14)) xor (A(93) and B(13)) xor (A(94) and B(12)) xor (A(95) and B(11)) xor (A(96) and B(10)) xor (A(97) and B(9)) xor (A(98) and B(8)) xor (A(99) and B(7)) xor (A(100) and B(6)) xor (A(101) and B(5)) xor (A(102) and B(4)) xor (A(103) and B(3)) xor (A(104) and B(2)) xor (A(105) and B(1)) xor (A(106) and B(0)) xor (A(99) and B(127)) xor (A(100) and B(126)) xor (A(101) and B(125)) xor (A(102) and B(124)) xor (A(103) and B(123)) xor (A(104) and B(122)) xor (A(105) and B(121)) xor (A(106) and B(120)) xor (A(107) and B(119)) xor (A(108) and B(118)) xor (A(109) and B(117)) xor (A(110) and B(116)) xor (A(111) and B(115)) xor (A(112) and B(114)) xor (A(113) and B(113)) xor (A(114) and B(112)) xor (A(115) and B(111)) xor (A(116) and B(110)) xor (A(117) and B(109)) xor (A(118) and B(108)) xor (A(119) and B(107)) xor (A(120) and B(106)) xor (A(121) and B(105)) xor (A(122) and B(104)) xor (A(123) and B(103)) xor (A(124) and B(102)) xor (A(125) and B(101)) xor (A(126) and B(100)) xor (A(104) and B(127)) xor (A(105) and B(126)) xor (A(106) and B(125)) xor (A(107) and B(124)) xor (A(108) and B(123)) xor (A(109) and B(122)) xor (A(110) and B(121)) xor (A(111) and B(120)) xor (A(112) and B(119)) xor (A(113) and B(118)) xor (A(114) and B(117)) xor (A(115) and B(116)) xor (A(116) and B(115)) xor (A(117) and B(114)) xor (A(118) and B(113)) xor (A(119) and B(112)) xor (A(120) and B(111)) xor (A(121) and B(110)) xor (A(122) and B(109)) xor (A(123) and B(108)) xor (A(124) and B(107)) xor (A(125) and B(106)) xor (A(126) and B(105)) xor (A(105) and B(127)) xor (A(106) and B(126)) xor (A(107) and B(125)) xor (A(108) and B(124)) xor (A(109) and B(123)) xor (A(110) and B(122)) xor (A(111) and B(121)) xor (A(112) and B(120)) xor (A(113) and B(119)) xor (A(114) and B(118)) xor (A(115) and B(117)) xor (A(116) and B(116)) xor (A(117) and B(115)) xor (A(118) and B(114)) xor (A(119) and B(113)) xor (A(120) and B(112)) xor (A(121) and B(111)) xor (A(122) and B(110)) xor (A(123) and B(109)) xor (A(124) and B(108)) xor (A(125) and B(107)) xor (A(126) and B(106)) xor (A(106) and B(127)) xor (A(107) and B(126)) xor (A(108) and B(125)) xor (A(109) and B(124)) xor (A(110) and B(123)) xor (A(111) and B(122)) xor (A(112) and B(121)) xor (A(113) and B(120)) xor (A(114) and B(119)) xor (A(115) and B(118)) xor (A(116) and B(117)) xor (A(117) and B(116)) xor (A(118) and B(115)) xor (A(119) and B(114)) xor (A(120) and B(113)) xor (A(121) and B(112)) xor (A(122) and B(111)) xor (A(123) and B(110)) xor (A(124) and B(109)) xor (A(125) and B(108)) xor (A(126) and B(108));
    C(107) <= (A(0) and B(107)) xor (A(1) and B(106)) xor (A(2) and B(105)) xor (A(3) and B(104)) xor (A(4) and B(103)) xor (A(5) and B(102)) xor (A(6) and B(101)) xor (A(7) and B(100)) xor (A(8) and B(99)) xor (A(9) and B(98)) xor (A(10) and B(97)) xor (A(11) and B(96)) xor (A(12) and B(95)) xor (A(13) and B(94)) xor (A(14) and B(93)) xor (A(15) and B(92)) xor (A(16) and B(91)) xor (A(17) and B(90)) xor (A(18) and B(89)) xor (A(19) and B(88)) xor (A(20) and B(87)) xor (A(21) and B(86)) xor (A(23) and B(85)) xor (A(23) and B(84)) xor (A(24) and B(83)) xor (A(25) and B(82)) xor (A(26) and B(81)) xor (A(27) and B(80)) xor (A(28) and B(79)) xor (A(29) and B(78)) xor (A(30) and B(77)) xor (A(31) and B(76)) xor (A(32) and B(75)) xor (A(33) and B(74)) xor (A(34) and B(73)) xor (A(35) and B(72)) xor (A(36) and B(71)) xor (A(37) and B(70)) xor (A(38) and B(69)) xor (A(39) and B(68)) xor (A(40) and B(67)) xor (A(41) and B(66)) xor (A(42) and B(65)) xor (A(43) and B(64)) xor (A(44) and B(63)) xor (A(45) and B(62)) xor (A(46) and B(61)) xor (A(47) and B(60)) xor (A(48) and B(59)) xor (A(49) and B(58)) xor (A(50) and B(57)) xor (A(51) and B(56)) xor (A(52) and B(55)) xor (A(53) and B(54)) xor (A(54) and B(53)) xor (A(55) and B(52)) xor (A(56) and B(51)) xor (A(57) and B(50)) xor (A(58) and B(49)) xor (A(59) and B(48)) xor (A(60) and B(47)) xor (A(61) and B(46)) xor (A(62) and B(45)) xor (A(63) and B(44)) xor (A(64) and B(43)) xor (A(65) and B(42)) xor (A(66) and B(41)) xor (A(67) and B(40)) xor (A(68) and B(39)) xor (A(69) and B(38)) xor (A(70) and B(37)) xor (A(71) and B(36)) xor (A(72) and B(35)) xor (A(73) and B(34)) xor (A(74) and B(33)) xor (A(75) and B(32)) xor (A(76) and B(31)) xor (A(77) and B(30)) xor (A(78) and B(29)) xor (A(79) and B(28)) xor (A(80) and B(27)) xor (A(81) and B(26)) xor (A(82) and B(25)) xor (A(83) and B(24)) xor (A(84) and B(23)) xor (A(85) and B(23)) xor (A(86) and B(21)) xor (A(87) and B(20)) xor (A(88) and B(19)) xor (A(89) and B(18)) xor (A(90) and B(17)) xor (A(91) and B(16)) xor (A(92) and B(15)) xor (A(93) and B(14)) xor (A(94) and B(13)) xor (A(95) and B(12)) xor (A(96) and B(11)) xor (A(97) and B(10)) xor (A(98) and B(9)) xor (A(99) and B(8)) xor (A(100) and B(7)) xor (A(101) and B(6)) xor (A(102) and B(5)) xor (A(103) and B(4)) xor (A(104) and B(3)) xor (A(105) and B(2)) xor (A(106) and B(1)) xor (A(107) and B(0)) xor (A(100) and B(127)) xor (A(101) and B(126)) xor (A(102) and B(125)) xor (A(103) and B(124)) xor (A(104) and B(123)) xor (A(105) and B(122)) xor (A(106) and B(121)) xor (A(107) and B(120)) xor (A(108) and B(119)) xor (A(109) and B(118)) xor (A(110) and B(117)) xor (A(111) and B(116)) xor (A(112) and B(115)) xor (A(113) and B(114)) xor (A(114) and B(113)) xor (A(115) and B(112)) xor (A(116) and B(111)) xor (A(117) and B(110)) xor (A(118) and B(109)) xor (A(119) and B(108)) xor (A(120) and B(107)) xor (A(121) and B(106)) xor (A(122) and B(105)) xor (A(123) and B(104)) xor (A(124) and B(103)) xor (A(125) and B(102)) xor (A(126) and B(101)) xor (A(105) and B(127)) xor (A(106) and B(126)) xor (A(107) and B(125)) xor (A(108) and B(124)) xor (A(109) and B(123)) xor (A(110) and B(122)) xor (A(111) and B(121)) xor (A(112) and B(120)) xor (A(113) and B(119)) xor (A(114) and B(118)) xor (A(115) and B(117)) xor (A(116) and B(116)) xor (A(117) and B(115)) xor (A(118) and B(114)) xor (A(119) and B(113)) xor (A(120) and B(112)) xor (A(121) and B(111)) xor (A(122) and B(110)) xor (A(123) and B(109)) xor (A(124) and B(108)) xor (A(125) and B(107)) xor (A(126) and B(106)) xor (A(106) and B(127)) xor (A(107) and B(126)) xor (A(108) and B(125)) xor (A(109) and B(124)) xor (A(110) and B(123)) xor (A(111) and B(122)) xor (A(112) and B(121)) xor (A(113) and B(120)) xor (A(114) and B(119)) xor (A(115) and B(118)) xor (A(116) and B(117)) xor (A(117) and B(116)) xor (A(118) and B(115)) xor (A(119) and B(114)) xor (A(120) and B(113)) xor (A(121) and B(112)) xor (A(122) and B(111)) xor (A(123) and B(110)) xor (A(124) and B(109)) xor (A(125) and B(108)) xor (A(126) and B(107)) xor (A(107) and B(127)) xor (A(108) and B(126)) xor (A(109) and B(125)) xor (A(110) and B(124)) xor (A(111) and B(123)) xor (A(112) and B(122)) xor (A(113) and B(121)) xor (A(114) and B(120)) xor (A(115) and B(119)) xor (A(116) and B(118)) xor (A(117) and B(117)) xor (A(118) and B(116)) xor (A(119) and B(115)) xor (A(120) and B(114)) xor (A(121) and B(113)) xor (A(122) and B(112)) xor (A(123) and B(111)) xor (A(124) and B(110)) xor (A(125) and B(109)) xor (A(126) and B(109));
    C(108) <= (A(0) and B(108)) xor (A(1) and B(107)) xor (A(2) and B(106)) xor (A(3) and B(105)) xor (A(4) and B(104)) xor (A(5) and B(103)) xor (A(6) and B(102)) xor (A(7) and B(101)) xor (A(8) and B(100)) xor (A(9) and B(99)) xor (A(10) and B(98)) xor (A(11) and B(97)) xor (A(12) and B(96)) xor (A(13) and B(95)) xor (A(14) and B(94)) xor (A(15) and B(93)) xor (A(16) and B(92)) xor (A(17) and B(91)) xor (A(18) and B(90)) xor (A(19) and B(89)) xor (A(20) and B(88)) xor (A(21) and B(87)) xor (A(23) and B(86)) xor (A(23) and B(85)) xor (A(24) and B(84)) xor (A(25) and B(83)) xor (A(26) and B(82)) xor (A(27) and B(81)) xor (A(28) and B(80)) xor (A(29) and B(79)) xor (A(30) and B(78)) xor (A(31) and B(77)) xor (A(32) and B(76)) xor (A(33) and B(75)) xor (A(34) and B(74)) xor (A(35) and B(73)) xor (A(36) and B(72)) xor (A(37) and B(71)) xor (A(38) and B(70)) xor (A(39) and B(69)) xor (A(40) and B(68)) xor (A(41) and B(67)) xor (A(42) and B(66)) xor (A(43) and B(65)) xor (A(44) and B(64)) xor (A(45) and B(63)) xor (A(46) and B(62)) xor (A(47) and B(61)) xor (A(48) and B(60)) xor (A(49) and B(59)) xor (A(50) and B(58)) xor (A(51) and B(57)) xor (A(52) and B(56)) xor (A(53) and B(55)) xor (A(54) and B(54)) xor (A(55) and B(53)) xor (A(56) and B(52)) xor (A(57) and B(51)) xor (A(58) and B(50)) xor (A(59) and B(49)) xor (A(60) and B(48)) xor (A(61) and B(47)) xor (A(62) and B(46)) xor (A(63) and B(45)) xor (A(64) and B(44)) xor (A(65) and B(43)) xor (A(66) and B(42)) xor (A(67) and B(41)) xor (A(68) and B(40)) xor (A(69) and B(39)) xor (A(70) and B(38)) xor (A(71) and B(37)) xor (A(72) and B(36)) xor (A(73) and B(35)) xor (A(74) and B(34)) xor (A(75) and B(33)) xor (A(76) and B(32)) xor (A(77) and B(31)) xor (A(78) and B(30)) xor (A(79) and B(29)) xor (A(80) and B(28)) xor (A(81) and B(27)) xor (A(82) and B(26)) xor (A(83) and B(25)) xor (A(84) and B(24)) xor (A(85) and B(23)) xor (A(86) and B(23)) xor (A(87) and B(21)) xor (A(88) and B(20)) xor (A(89) and B(19)) xor (A(90) and B(18)) xor (A(91) and B(17)) xor (A(92) and B(16)) xor (A(93) and B(15)) xor (A(94) and B(14)) xor (A(95) and B(13)) xor (A(96) and B(12)) xor (A(97) and B(11)) xor (A(98) and B(10)) xor (A(99) and B(9)) xor (A(100) and B(8)) xor (A(101) and B(7)) xor (A(102) and B(6)) xor (A(103) and B(5)) xor (A(104) and B(4)) xor (A(105) and B(3)) xor (A(106) and B(2)) xor (A(107) and B(1)) xor (A(108) and B(0)) xor (A(101) and B(127)) xor (A(102) and B(126)) xor (A(103) and B(125)) xor (A(104) and B(124)) xor (A(105) and B(123)) xor (A(106) and B(122)) xor (A(107) and B(121)) xor (A(108) and B(120)) xor (A(109) and B(119)) xor (A(110) and B(118)) xor (A(111) and B(117)) xor (A(112) and B(116)) xor (A(113) and B(115)) xor (A(114) and B(114)) xor (A(115) and B(113)) xor (A(116) and B(112)) xor (A(117) and B(111)) xor (A(118) and B(110)) xor (A(119) and B(109)) xor (A(120) and B(108)) xor (A(121) and B(107)) xor (A(122) and B(106)) xor (A(123) and B(105)) xor (A(124) and B(104)) xor (A(125) and B(103)) xor (A(126) and B(102)) xor (A(106) and B(127)) xor (A(107) and B(126)) xor (A(108) and B(125)) xor (A(109) and B(124)) xor (A(110) and B(123)) xor (A(111) and B(122)) xor (A(112) and B(121)) xor (A(113) and B(120)) xor (A(114) and B(119)) xor (A(115) and B(118)) xor (A(116) and B(117)) xor (A(117) and B(116)) xor (A(118) and B(115)) xor (A(119) and B(114)) xor (A(120) and B(113)) xor (A(121) and B(112)) xor (A(122) and B(111)) xor (A(123) and B(110)) xor (A(124) and B(109)) xor (A(125) and B(108)) xor (A(126) and B(107)) xor (A(107) and B(127)) xor (A(108) and B(126)) xor (A(109) and B(125)) xor (A(110) and B(124)) xor (A(111) and B(123)) xor (A(112) and B(122)) xor (A(113) and B(121)) xor (A(114) and B(120)) xor (A(115) and B(119)) xor (A(116) and B(118)) xor (A(117) and B(117)) xor (A(118) and B(116)) xor (A(119) and B(115)) xor (A(120) and B(114)) xor (A(121) and B(113)) xor (A(122) and B(112)) xor (A(123) and B(111)) xor (A(124) and B(110)) xor (A(125) and B(109)) xor (A(126) and B(108)) xor (A(108) and B(127)) xor (A(109) and B(126)) xor (A(110) and B(125)) xor (A(111) and B(124)) xor (A(112) and B(123)) xor (A(113) and B(122)) xor (A(114) and B(121)) xor (A(115) and B(120)) xor (A(116) and B(119)) xor (A(117) and B(118)) xor (A(118) and B(117)) xor (A(119) and B(116)) xor (A(120) and B(115)) xor (A(121) and B(114)) xor (A(122) and B(113)) xor (A(123) and B(112)) xor (A(124) and B(111)) xor (A(125) and B(110)) xor (A(126) and B(110));
    C(109) <= (A(0) and B(109)) xor (A(1) and B(108)) xor (A(2) and B(107)) xor (A(3) and B(106)) xor (A(4) and B(105)) xor (A(5) and B(104)) xor (A(6) and B(103)) xor (A(7) and B(102)) xor (A(8) and B(101)) xor (A(9) and B(100)) xor (A(10) and B(99)) xor (A(11) and B(98)) xor (A(12) and B(97)) xor (A(13) and B(96)) xor (A(14) and B(95)) xor (A(15) and B(94)) xor (A(16) and B(93)) xor (A(17) and B(92)) xor (A(18) and B(91)) xor (A(19) and B(90)) xor (A(20) and B(89)) xor (A(21) and B(88)) xor (A(23) and B(87)) xor (A(23) and B(86)) xor (A(24) and B(85)) xor (A(25) and B(84)) xor (A(26) and B(83)) xor (A(27) and B(82)) xor (A(28) and B(81)) xor (A(29) and B(80)) xor (A(30) and B(79)) xor (A(31) and B(78)) xor (A(32) and B(77)) xor (A(33) and B(76)) xor (A(34) and B(75)) xor (A(35) and B(74)) xor (A(36) and B(73)) xor (A(37) and B(72)) xor (A(38) and B(71)) xor (A(39) and B(70)) xor (A(40) and B(69)) xor (A(41) and B(68)) xor (A(42) and B(67)) xor (A(43) and B(66)) xor (A(44) and B(65)) xor (A(45) and B(64)) xor (A(46) and B(63)) xor (A(47) and B(62)) xor (A(48) and B(61)) xor (A(49) and B(60)) xor (A(50) and B(59)) xor (A(51) and B(58)) xor (A(52) and B(57)) xor (A(53) and B(56)) xor (A(54) and B(55)) xor (A(55) and B(54)) xor (A(56) and B(53)) xor (A(57) and B(52)) xor (A(58) and B(51)) xor (A(59) and B(50)) xor (A(60) and B(49)) xor (A(61) and B(48)) xor (A(62) and B(47)) xor (A(63) and B(46)) xor (A(64) and B(45)) xor (A(65) and B(44)) xor (A(66) and B(43)) xor (A(67) and B(42)) xor (A(68) and B(41)) xor (A(69) and B(40)) xor (A(70) and B(39)) xor (A(71) and B(38)) xor (A(72) and B(37)) xor (A(73) and B(36)) xor (A(74) and B(35)) xor (A(75) and B(34)) xor (A(76) and B(33)) xor (A(77) and B(32)) xor (A(78) and B(31)) xor (A(79) and B(30)) xor (A(80) and B(29)) xor (A(81) and B(28)) xor (A(82) and B(27)) xor (A(83) and B(26)) xor (A(84) and B(25)) xor (A(85) and B(24)) xor (A(86) and B(23)) xor (A(87) and B(23)) xor (A(88) and B(21)) xor (A(89) and B(20)) xor (A(90) and B(19)) xor (A(91) and B(18)) xor (A(92) and B(17)) xor (A(93) and B(16)) xor (A(94) and B(15)) xor (A(95) and B(14)) xor (A(96) and B(13)) xor (A(97) and B(12)) xor (A(98) and B(11)) xor (A(99) and B(10)) xor (A(100) and B(9)) xor (A(101) and B(8)) xor (A(102) and B(7)) xor (A(103) and B(6)) xor (A(104) and B(5)) xor (A(105) and B(4)) xor (A(106) and B(3)) xor (A(107) and B(2)) xor (A(108) and B(1)) xor (A(109) and B(0)) xor (A(102) and B(127)) xor (A(103) and B(126)) xor (A(104) and B(125)) xor (A(105) and B(124)) xor (A(106) and B(123)) xor (A(107) and B(122)) xor (A(108) and B(121)) xor (A(109) and B(120)) xor (A(110) and B(119)) xor (A(111) and B(118)) xor (A(112) and B(117)) xor (A(113) and B(116)) xor (A(114) and B(115)) xor (A(115) and B(114)) xor (A(116) and B(113)) xor (A(117) and B(112)) xor (A(118) and B(111)) xor (A(119) and B(110)) xor (A(120) and B(109)) xor (A(121) and B(108)) xor (A(122) and B(107)) xor (A(123) and B(106)) xor (A(124) and B(105)) xor (A(125) and B(104)) xor (A(126) and B(103)) xor (A(107) and B(127)) xor (A(108) and B(126)) xor (A(109) and B(125)) xor (A(110) and B(124)) xor (A(111) and B(123)) xor (A(112) and B(122)) xor (A(113) and B(121)) xor (A(114) and B(120)) xor (A(115) and B(119)) xor (A(116) and B(118)) xor (A(117) and B(117)) xor (A(118) and B(116)) xor (A(119) and B(115)) xor (A(120) and B(114)) xor (A(121) and B(113)) xor (A(122) and B(112)) xor (A(123) and B(111)) xor (A(124) and B(110)) xor (A(125) and B(109)) xor (A(126) and B(108)) xor (A(108) and B(127)) xor (A(109) and B(126)) xor (A(110) and B(125)) xor (A(111) and B(124)) xor (A(112) and B(123)) xor (A(113) and B(122)) xor (A(114) and B(121)) xor (A(115) and B(120)) xor (A(116) and B(119)) xor (A(117) and B(118)) xor (A(118) and B(117)) xor (A(119) and B(116)) xor (A(120) and B(115)) xor (A(121) and B(114)) xor (A(122) and B(113)) xor (A(123) and B(112)) xor (A(124) and B(111)) xor (A(125) and B(110)) xor (A(126) and B(109)) xor (A(109) and B(127)) xor (A(110) and B(126)) xor (A(111) and B(125)) xor (A(112) and B(124)) xor (A(113) and B(123)) xor (A(114) and B(122)) xor (A(115) and B(121)) xor (A(116) and B(120)) xor (A(117) and B(119)) xor (A(118) and B(118)) xor (A(119) and B(117)) xor (A(120) and B(116)) xor (A(121) and B(115)) xor (A(122) and B(114)) xor (A(123) and B(113)) xor (A(124) and B(112)) xor (A(125) and B(111)) xor (A(126) and B(111));
    C(110) <= (A(0) and B(110)) xor (A(1) and B(109)) xor (A(2) and B(108)) xor (A(3) and B(107)) xor (A(4) and B(106)) xor (A(5) and B(105)) xor (A(6) and B(104)) xor (A(7) and B(103)) xor (A(8) and B(102)) xor (A(9) and B(101)) xor (A(10) and B(100)) xor (A(11) and B(99)) xor (A(12) and B(98)) xor (A(13) and B(97)) xor (A(14) and B(96)) xor (A(15) and B(95)) xor (A(16) and B(94)) xor (A(17) and B(93)) xor (A(18) and B(92)) xor (A(19) and B(91)) xor (A(20) and B(90)) xor (A(21) and B(89)) xor (A(23) and B(88)) xor (A(23) and B(87)) xor (A(24) and B(86)) xor (A(25) and B(85)) xor (A(26) and B(84)) xor (A(27) and B(83)) xor (A(28) and B(82)) xor (A(29) and B(81)) xor (A(30) and B(80)) xor (A(31) and B(79)) xor (A(32) and B(78)) xor (A(33) and B(77)) xor (A(34) and B(76)) xor (A(35) and B(75)) xor (A(36) and B(74)) xor (A(37) and B(73)) xor (A(38) and B(72)) xor (A(39) and B(71)) xor (A(40) and B(70)) xor (A(41) and B(69)) xor (A(42) and B(68)) xor (A(43) and B(67)) xor (A(44) and B(66)) xor (A(45) and B(65)) xor (A(46) and B(64)) xor (A(47) and B(63)) xor (A(48) and B(62)) xor (A(49) and B(61)) xor (A(50) and B(60)) xor (A(51) and B(59)) xor (A(52) and B(58)) xor (A(53) and B(57)) xor (A(54) and B(56)) xor (A(55) and B(55)) xor (A(56) and B(54)) xor (A(57) and B(53)) xor (A(58) and B(52)) xor (A(59) and B(51)) xor (A(60) and B(50)) xor (A(61) and B(49)) xor (A(62) and B(48)) xor (A(63) and B(47)) xor (A(64) and B(46)) xor (A(65) and B(45)) xor (A(66) and B(44)) xor (A(67) and B(43)) xor (A(68) and B(42)) xor (A(69) and B(41)) xor (A(70) and B(40)) xor (A(71) and B(39)) xor (A(72) and B(38)) xor (A(73) and B(37)) xor (A(74) and B(36)) xor (A(75) and B(35)) xor (A(76) and B(34)) xor (A(77) and B(33)) xor (A(78) and B(32)) xor (A(79) and B(31)) xor (A(80) and B(30)) xor (A(81) and B(29)) xor (A(82) and B(28)) xor (A(83) and B(27)) xor (A(84) and B(26)) xor (A(85) and B(25)) xor (A(86) and B(24)) xor (A(87) and B(23)) xor (A(88) and B(23)) xor (A(89) and B(21)) xor (A(90) and B(20)) xor (A(91) and B(19)) xor (A(92) and B(18)) xor (A(93) and B(17)) xor (A(94) and B(16)) xor (A(95) and B(15)) xor (A(96) and B(14)) xor (A(97) and B(13)) xor (A(98) and B(12)) xor (A(99) and B(11)) xor (A(100) and B(10)) xor (A(101) and B(9)) xor (A(102) and B(8)) xor (A(103) and B(7)) xor (A(104) and B(6)) xor (A(105) and B(5)) xor (A(106) and B(4)) xor (A(107) and B(3)) xor (A(108) and B(2)) xor (A(109) and B(1)) xor (A(110) and B(0)) xor (A(103) and B(127)) xor (A(104) and B(126)) xor (A(105) and B(125)) xor (A(106) and B(124)) xor (A(107) and B(123)) xor (A(108) and B(122)) xor (A(109) and B(121)) xor (A(110) and B(120)) xor (A(111) and B(119)) xor (A(112) and B(118)) xor (A(113) and B(117)) xor (A(114) and B(116)) xor (A(115) and B(115)) xor (A(116) and B(114)) xor (A(117) and B(113)) xor (A(118) and B(112)) xor (A(119) and B(111)) xor (A(120) and B(110)) xor (A(121) and B(109)) xor (A(122) and B(108)) xor (A(123) and B(107)) xor (A(124) and B(106)) xor (A(125) and B(105)) xor (A(126) and B(104)) xor (A(108) and B(127)) xor (A(109) and B(126)) xor (A(110) and B(125)) xor (A(111) and B(124)) xor (A(112) and B(123)) xor (A(113) and B(122)) xor (A(114) and B(121)) xor (A(115) and B(120)) xor (A(116) and B(119)) xor (A(117) and B(118)) xor (A(118) and B(117)) xor (A(119) and B(116)) xor (A(120) and B(115)) xor (A(121) and B(114)) xor (A(122) and B(113)) xor (A(123) and B(112)) xor (A(124) and B(111)) xor (A(125) and B(110)) xor (A(126) and B(109)) xor (A(109) and B(127)) xor (A(110) and B(126)) xor (A(111) and B(125)) xor (A(112) and B(124)) xor (A(113) and B(123)) xor (A(114) and B(122)) xor (A(115) and B(121)) xor (A(116) and B(120)) xor (A(117) and B(119)) xor (A(118) and B(118)) xor (A(119) and B(117)) xor (A(120) and B(116)) xor (A(121) and B(115)) xor (A(122) and B(114)) xor (A(123) and B(113)) xor (A(124) and B(112)) xor (A(125) and B(111)) xor (A(126) and B(110)) xor (A(110) and B(127)) xor (A(111) and B(126)) xor (A(112) and B(125)) xor (A(113) and B(124)) xor (A(114) and B(123)) xor (A(115) and B(122)) xor (A(116) and B(121)) xor (A(117) and B(120)) xor (A(118) and B(119)) xor (A(119) and B(118)) xor (A(120) and B(117)) xor (A(121) and B(116)) xor (A(122) and B(115)) xor (A(123) and B(114)) xor (A(124) and B(113)) xor (A(125) and B(112)) xor (A(126) and B(112));
    C(111) <= (A(0) and B(111)) xor (A(1) and B(110)) xor (A(2) and B(109)) xor (A(3) and B(108)) xor (A(4) and B(107)) xor (A(5) and B(106)) xor (A(6) and B(105)) xor (A(7) and B(104)) xor (A(8) and B(103)) xor (A(9) and B(102)) xor (A(10) and B(101)) xor (A(11) and B(100)) xor (A(12) and B(99)) xor (A(13) and B(98)) xor (A(14) and B(97)) xor (A(15) and B(96)) xor (A(16) and B(95)) xor (A(17) and B(94)) xor (A(18) and B(93)) xor (A(19) and B(92)) xor (A(20) and B(91)) xor (A(21) and B(90)) xor (A(23) and B(89)) xor (A(23) and B(88)) xor (A(24) and B(87)) xor (A(25) and B(86)) xor (A(26) and B(85)) xor (A(27) and B(84)) xor (A(28) and B(83)) xor (A(29) and B(82)) xor (A(30) and B(81)) xor (A(31) and B(80)) xor (A(32) and B(79)) xor (A(33) and B(78)) xor (A(34) and B(77)) xor (A(35) and B(76)) xor (A(36) and B(75)) xor (A(37) and B(74)) xor (A(38) and B(73)) xor (A(39) and B(72)) xor (A(40) and B(71)) xor (A(41) and B(70)) xor (A(42) and B(69)) xor (A(43) and B(68)) xor (A(44) and B(67)) xor (A(45) and B(66)) xor (A(46) and B(65)) xor (A(47) and B(64)) xor (A(48) and B(63)) xor (A(49) and B(62)) xor (A(50) and B(61)) xor (A(51) and B(60)) xor (A(52) and B(59)) xor (A(53) and B(58)) xor (A(54) and B(57)) xor (A(55) and B(56)) xor (A(56) and B(55)) xor (A(57) and B(54)) xor (A(58) and B(53)) xor (A(59) and B(52)) xor (A(60) and B(51)) xor (A(61) and B(50)) xor (A(62) and B(49)) xor (A(63) and B(48)) xor (A(64) and B(47)) xor (A(65) and B(46)) xor (A(66) and B(45)) xor (A(67) and B(44)) xor (A(68) and B(43)) xor (A(69) and B(42)) xor (A(70) and B(41)) xor (A(71) and B(40)) xor (A(72) and B(39)) xor (A(73) and B(38)) xor (A(74) and B(37)) xor (A(75) and B(36)) xor (A(76) and B(35)) xor (A(77) and B(34)) xor (A(78) and B(33)) xor (A(79) and B(32)) xor (A(80) and B(31)) xor (A(81) and B(30)) xor (A(82) and B(29)) xor (A(83) and B(28)) xor (A(84) and B(27)) xor (A(85) and B(26)) xor (A(86) and B(25)) xor (A(87) and B(24)) xor (A(88) and B(23)) xor (A(89) and B(23)) xor (A(90) and B(21)) xor (A(91) and B(20)) xor (A(92) and B(19)) xor (A(93) and B(18)) xor (A(94) and B(17)) xor (A(95) and B(16)) xor (A(96) and B(15)) xor (A(97) and B(14)) xor (A(98) and B(13)) xor (A(99) and B(12)) xor (A(100) and B(11)) xor (A(101) and B(10)) xor (A(102) and B(9)) xor (A(103) and B(8)) xor (A(104) and B(7)) xor (A(105) and B(6)) xor (A(106) and B(5)) xor (A(107) and B(4)) xor (A(108) and B(3)) xor (A(109) and B(2)) xor (A(110) and B(1)) xor (A(111) and B(0)) xor (A(104) and B(127)) xor (A(105) and B(126)) xor (A(106) and B(125)) xor (A(107) and B(124)) xor (A(108) and B(123)) xor (A(109) and B(122)) xor (A(110) and B(121)) xor (A(111) and B(120)) xor (A(112) and B(119)) xor (A(113) and B(118)) xor (A(114) and B(117)) xor (A(115) and B(116)) xor (A(116) and B(115)) xor (A(117) and B(114)) xor (A(118) and B(113)) xor (A(119) and B(112)) xor (A(120) and B(111)) xor (A(121) and B(110)) xor (A(122) and B(109)) xor (A(123) and B(108)) xor (A(124) and B(107)) xor (A(125) and B(106)) xor (A(126) and B(105)) xor (A(109) and B(127)) xor (A(110) and B(126)) xor (A(111) and B(125)) xor (A(112) and B(124)) xor (A(113) and B(123)) xor (A(114) and B(122)) xor (A(115) and B(121)) xor (A(116) and B(120)) xor (A(117) and B(119)) xor (A(118) and B(118)) xor (A(119) and B(117)) xor (A(120) and B(116)) xor (A(121) and B(115)) xor (A(122) and B(114)) xor (A(123) and B(113)) xor (A(124) and B(112)) xor (A(125) and B(111)) xor (A(126) and B(110)) xor (A(110) and B(127)) xor (A(111) and B(126)) xor (A(112) and B(125)) xor (A(113) and B(124)) xor (A(114) and B(123)) xor (A(115) and B(122)) xor (A(116) and B(121)) xor (A(117) and B(120)) xor (A(118) and B(119)) xor (A(119) and B(118)) xor (A(120) and B(117)) xor (A(121) and B(116)) xor (A(122) and B(115)) xor (A(123) and B(114)) xor (A(124) and B(113)) xor (A(125) and B(112)) xor (A(126) and B(111)) xor (A(111) and B(127)) xor (A(112) and B(126)) xor (A(113) and B(125)) xor (A(114) and B(124)) xor (A(115) and B(123)) xor (A(116) and B(122)) xor (A(117) and B(121)) xor (A(118) and B(120)) xor (A(119) and B(119)) xor (A(120) and B(118)) xor (A(121) and B(117)) xor (A(122) and B(116)) xor (A(123) and B(115)) xor (A(124) and B(114)) xor (A(125) and B(113)) xor (A(126) and B(113));
    C(112) <= (A(0) and B(112)) xor (A(1) and B(111)) xor (A(2) and B(110)) xor (A(3) and B(109)) xor (A(4) and B(108)) xor (A(5) and B(107)) xor (A(6) and B(106)) xor (A(7) and B(105)) xor (A(8) and B(104)) xor (A(9) and B(103)) xor (A(10) and B(102)) xor (A(11) and B(101)) xor (A(12) and B(100)) xor (A(13) and B(99)) xor (A(14) and B(98)) xor (A(15) and B(97)) xor (A(16) and B(96)) xor (A(17) and B(95)) xor (A(18) and B(94)) xor (A(19) and B(93)) xor (A(20) and B(92)) xor (A(21) and B(91)) xor (A(23) and B(90)) xor (A(23) and B(89)) xor (A(24) and B(88)) xor (A(25) and B(87)) xor (A(26) and B(86)) xor (A(27) and B(85)) xor (A(28) and B(84)) xor (A(29) and B(83)) xor (A(30) and B(82)) xor (A(31) and B(81)) xor (A(32) and B(80)) xor (A(33) and B(79)) xor (A(34) and B(78)) xor (A(35) and B(77)) xor (A(36) and B(76)) xor (A(37) and B(75)) xor (A(38) and B(74)) xor (A(39) and B(73)) xor (A(40) and B(72)) xor (A(41) and B(71)) xor (A(42) and B(70)) xor (A(43) and B(69)) xor (A(44) and B(68)) xor (A(45) and B(67)) xor (A(46) and B(66)) xor (A(47) and B(65)) xor (A(48) and B(64)) xor (A(49) and B(63)) xor (A(50) and B(62)) xor (A(51) and B(61)) xor (A(52) and B(60)) xor (A(53) and B(59)) xor (A(54) and B(58)) xor (A(55) and B(57)) xor (A(56) and B(56)) xor (A(57) and B(55)) xor (A(58) and B(54)) xor (A(59) and B(53)) xor (A(60) and B(52)) xor (A(61) and B(51)) xor (A(62) and B(50)) xor (A(63) and B(49)) xor (A(64) and B(48)) xor (A(65) and B(47)) xor (A(66) and B(46)) xor (A(67) and B(45)) xor (A(68) and B(44)) xor (A(69) and B(43)) xor (A(70) and B(42)) xor (A(71) and B(41)) xor (A(72) and B(40)) xor (A(73) and B(39)) xor (A(74) and B(38)) xor (A(75) and B(37)) xor (A(76) and B(36)) xor (A(77) and B(35)) xor (A(78) and B(34)) xor (A(79) and B(33)) xor (A(80) and B(32)) xor (A(81) and B(31)) xor (A(82) and B(30)) xor (A(83) and B(29)) xor (A(84) and B(28)) xor (A(85) and B(27)) xor (A(86) and B(26)) xor (A(87) and B(25)) xor (A(88) and B(24)) xor (A(89) and B(23)) xor (A(90) and B(23)) xor (A(91) and B(21)) xor (A(92) and B(20)) xor (A(93) and B(19)) xor (A(94) and B(18)) xor (A(95) and B(17)) xor (A(96) and B(16)) xor (A(97) and B(15)) xor (A(98) and B(14)) xor (A(99) and B(13)) xor (A(100) and B(12)) xor (A(101) and B(11)) xor (A(102) and B(10)) xor (A(103) and B(9)) xor (A(104) and B(8)) xor (A(105) and B(7)) xor (A(106) and B(6)) xor (A(107) and B(5)) xor (A(108) and B(4)) xor (A(109) and B(3)) xor (A(110) and B(2)) xor (A(111) and B(1)) xor (A(112) and B(0)) xor (A(105) and B(127)) xor (A(106) and B(126)) xor (A(107) and B(125)) xor (A(108) and B(124)) xor (A(109) and B(123)) xor (A(110) and B(122)) xor (A(111) and B(121)) xor (A(112) and B(120)) xor (A(113) and B(119)) xor (A(114) and B(118)) xor (A(115) and B(117)) xor (A(116) and B(116)) xor (A(117) and B(115)) xor (A(118) and B(114)) xor (A(119) and B(113)) xor (A(120) and B(112)) xor (A(121) and B(111)) xor (A(122) and B(110)) xor (A(123) and B(109)) xor (A(124) and B(108)) xor (A(125) and B(107)) xor (A(126) and B(106)) xor (A(110) and B(127)) xor (A(111) and B(126)) xor (A(112) and B(125)) xor (A(113) and B(124)) xor (A(114) and B(123)) xor (A(115) and B(122)) xor (A(116) and B(121)) xor (A(117) and B(120)) xor (A(118) and B(119)) xor (A(119) and B(118)) xor (A(120) and B(117)) xor (A(121) and B(116)) xor (A(122) and B(115)) xor (A(123) and B(114)) xor (A(124) and B(113)) xor (A(125) and B(112)) xor (A(126) and B(111)) xor (A(111) and B(127)) xor (A(112) and B(126)) xor (A(113) and B(125)) xor (A(114) and B(124)) xor (A(115) and B(123)) xor (A(116) and B(122)) xor (A(117) and B(121)) xor (A(118) and B(120)) xor (A(119) and B(119)) xor (A(120) and B(118)) xor (A(121) and B(117)) xor (A(122) and B(116)) xor (A(123) and B(115)) xor (A(124) and B(114)) xor (A(125) and B(113)) xor (A(126) and B(112)) xor (A(112) and B(127)) xor (A(113) and B(126)) xor (A(114) and B(125)) xor (A(115) and B(124)) xor (A(116) and B(123)) xor (A(117) and B(122)) xor (A(118) and B(121)) xor (A(119) and B(120)) xor (A(120) and B(119)) xor (A(121) and B(118)) xor (A(122) and B(117)) xor (A(123) and B(116)) xor (A(124) and B(115)) xor (A(125) and B(114)) xor (A(126) and B(114));
    C(113) <= (A(0) and B(113)) xor (A(1) and B(112)) xor (A(2) and B(111)) xor (A(3) and B(110)) xor (A(4) and B(109)) xor (A(5) and B(108)) xor (A(6) and B(107)) xor (A(7) and B(106)) xor (A(8) and B(105)) xor (A(9) and B(104)) xor (A(10) and B(103)) xor (A(11) and B(102)) xor (A(12) and B(101)) xor (A(13) and B(100)) xor (A(14) and B(99)) xor (A(15) and B(98)) xor (A(16) and B(97)) xor (A(17) and B(96)) xor (A(18) and B(95)) xor (A(19) and B(94)) xor (A(20) and B(93)) xor (A(21) and B(92)) xor (A(23) and B(91)) xor (A(23) and B(90)) xor (A(24) and B(89)) xor (A(25) and B(88)) xor (A(26) and B(87)) xor (A(27) and B(86)) xor (A(28) and B(85)) xor (A(29) and B(84)) xor (A(30) and B(83)) xor (A(31) and B(82)) xor (A(32) and B(81)) xor (A(33) and B(80)) xor (A(34) and B(79)) xor (A(35) and B(78)) xor (A(36) and B(77)) xor (A(37) and B(76)) xor (A(38) and B(75)) xor (A(39) and B(74)) xor (A(40) and B(73)) xor (A(41) and B(72)) xor (A(42) and B(71)) xor (A(43) and B(70)) xor (A(44) and B(69)) xor (A(45) and B(68)) xor (A(46) and B(67)) xor (A(47) and B(66)) xor (A(48) and B(65)) xor (A(49) and B(64)) xor (A(50) and B(63)) xor (A(51) and B(62)) xor (A(52) and B(61)) xor (A(53) and B(60)) xor (A(54) and B(59)) xor (A(55) and B(58)) xor (A(56) and B(57)) xor (A(57) and B(56)) xor (A(58) and B(55)) xor (A(59) and B(54)) xor (A(60) and B(53)) xor (A(61) and B(52)) xor (A(62) and B(51)) xor (A(63) and B(50)) xor (A(64) and B(49)) xor (A(65) and B(48)) xor (A(66) and B(47)) xor (A(67) and B(46)) xor (A(68) and B(45)) xor (A(69) and B(44)) xor (A(70) and B(43)) xor (A(71) and B(42)) xor (A(72) and B(41)) xor (A(73) and B(40)) xor (A(74) and B(39)) xor (A(75) and B(38)) xor (A(76) and B(37)) xor (A(77) and B(36)) xor (A(78) and B(35)) xor (A(79) and B(34)) xor (A(80) and B(33)) xor (A(81) and B(32)) xor (A(82) and B(31)) xor (A(83) and B(30)) xor (A(84) and B(29)) xor (A(85) and B(28)) xor (A(86) and B(27)) xor (A(87) and B(26)) xor (A(88) and B(25)) xor (A(89) and B(24)) xor (A(90) and B(23)) xor (A(91) and B(23)) xor (A(92) and B(21)) xor (A(93) and B(20)) xor (A(94) and B(19)) xor (A(95) and B(18)) xor (A(96) and B(17)) xor (A(97) and B(16)) xor (A(98) and B(15)) xor (A(99) and B(14)) xor (A(100) and B(13)) xor (A(101) and B(12)) xor (A(102) and B(11)) xor (A(103) and B(10)) xor (A(104) and B(9)) xor (A(105) and B(8)) xor (A(106) and B(7)) xor (A(107) and B(6)) xor (A(108) and B(5)) xor (A(109) and B(4)) xor (A(110) and B(3)) xor (A(111) and B(2)) xor (A(112) and B(1)) xor (A(113) and B(0)) xor (A(106) and B(127)) xor (A(107) and B(126)) xor (A(108) and B(125)) xor (A(109) and B(124)) xor (A(110) and B(123)) xor (A(111) and B(122)) xor (A(112) and B(121)) xor (A(113) and B(120)) xor (A(114) and B(119)) xor (A(115) and B(118)) xor (A(116) and B(117)) xor (A(117) and B(116)) xor (A(118) and B(115)) xor (A(119) and B(114)) xor (A(120) and B(113)) xor (A(121) and B(112)) xor (A(122) and B(111)) xor (A(123) and B(110)) xor (A(124) and B(109)) xor (A(125) and B(108)) xor (A(126) and B(107)) xor (A(111) and B(127)) xor (A(112) and B(126)) xor (A(113) and B(125)) xor (A(114) and B(124)) xor (A(115) and B(123)) xor (A(116) and B(122)) xor (A(117) and B(121)) xor (A(118) and B(120)) xor (A(119) and B(119)) xor (A(120) and B(118)) xor (A(121) and B(117)) xor (A(122) and B(116)) xor (A(123) and B(115)) xor (A(124) and B(114)) xor (A(125) and B(113)) xor (A(126) and B(112)) xor (A(112) and B(127)) xor (A(113) and B(126)) xor (A(114) and B(125)) xor (A(115) and B(124)) xor (A(116) and B(123)) xor (A(117) and B(122)) xor (A(118) and B(121)) xor (A(119) and B(120)) xor (A(120) and B(119)) xor (A(121) and B(118)) xor (A(122) and B(117)) xor (A(123) and B(116)) xor (A(124) and B(115)) xor (A(125) and B(114)) xor (A(126) and B(113)) xor (A(113) and B(127)) xor (A(114) and B(126)) xor (A(115) and B(125)) xor (A(116) and B(124)) xor (A(117) and B(123)) xor (A(118) and B(122)) xor (A(119) and B(121)) xor (A(120) and B(120)) xor (A(121) and B(119)) xor (A(122) and B(118)) xor (A(123) and B(117)) xor (A(124) and B(116)) xor (A(125) and B(115)) xor (A(126) and B(115));
    C(114) <= (A(0) and B(114)) xor (A(1) and B(113)) xor (A(2) and B(112)) xor (A(3) and B(111)) xor (A(4) and B(110)) xor (A(5) and B(109)) xor (A(6) and B(108)) xor (A(7) and B(107)) xor (A(8) and B(106)) xor (A(9) and B(105)) xor (A(10) and B(104)) xor (A(11) and B(103)) xor (A(12) and B(102)) xor (A(13) and B(101)) xor (A(14) and B(100)) xor (A(15) and B(99)) xor (A(16) and B(98)) xor (A(17) and B(97)) xor (A(18) and B(96)) xor (A(19) and B(95)) xor (A(20) and B(94)) xor (A(21) and B(93)) xor (A(23) and B(92)) xor (A(23) and B(91)) xor (A(24) and B(90)) xor (A(25) and B(89)) xor (A(26) and B(88)) xor (A(27) and B(87)) xor (A(28) and B(86)) xor (A(29) and B(85)) xor (A(30) and B(84)) xor (A(31) and B(83)) xor (A(32) and B(82)) xor (A(33) and B(81)) xor (A(34) and B(80)) xor (A(35) and B(79)) xor (A(36) and B(78)) xor (A(37) and B(77)) xor (A(38) and B(76)) xor (A(39) and B(75)) xor (A(40) and B(74)) xor (A(41) and B(73)) xor (A(42) and B(72)) xor (A(43) and B(71)) xor (A(44) and B(70)) xor (A(45) and B(69)) xor (A(46) and B(68)) xor (A(47) and B(67)) xor (A(48) and B(66)) xor (A(49) and B(65)) xor (A(50) and B(64)) xor (A(51) and B(63)) xor (A(52) and B(62)) xor (A(53) and B(61)) xor (A(54) and B(60)) xor (A(55) and B(59)) xor (A(56) and B(58)) xor (A(57) and B(57)) xor (A(58) and B(56)) xor (A(59) and B(55)) xor (A(60) and B(54)) xor (A(61) and B(53)) xor (A(62) and B(52)) xor (A(63) and B(51)) xor (A(64) and B(50)) xor (A(65) and B(49)) xor (A(66) and B(48)) xor (A(67) and B(47)) xor (A(68) and B(46)) xor (A(69) and B(45)) xor (A(70) and B(44)) xor (A(71) and B(43)) xor (A(72) and B(42)) xor (A(73) and B(41)) xor (A(74) and B(40)) xor (A(75) and B(39)) xor (A(76) and B(38)) xor (A(77) and B(37)) xor (A(78) and B(36)) xor (A(79) and B(35)) xor (A(80) and B(34)) xor (A(81) and B(33)) xor (A(82) and B(32)) xor (A(83) and B(31)) xor (A(84) and B(30)) xor (A(85) and B(29)) xor (A(86) and B(28)) xor (A(87) and B(27)) xor (A(88) and B(26)) xor (A(89) and B(25)) xor (A(90) and B(24)) xor (A(91) and B(23)) xor (A(92) and B(23)) xor (A(93) and B(21)) xor (A(94) and B(20)) xor (A(95) and B(19)) xor (A(96) and B(18)) xor (A(97) and B(17)) xor (A(98) and B(16)) xor (A(99) and B(15)) xor (A(100) and B(14)) xor (A(101) and B(13)) xor (A(102) and B(12)) xor (A(103) and B(11)) xor (A(104) and B(10)) xor (A(105) and B(9)) xor (A(106) and B(8)) xor (A(107) and B(7)) xor (A(108) and B(6)) xor (A(109) and B(5)) xor (A(110) and B(4)) xor (A(111) and B(3)) xor (A(112) and B(2)) xor (A(113) and B(1)) xor (A(114) and B(0)) xor (A(107) and B(127)) xor (A(108) and B(126)) xor (A(109) and B(125)) xor (A(110) and B(124)) xor (A(111) and B(123)) xor (A(112) and B(122)) xor (A(113) and B(121)) xor (A(114) and B(120)) xor (A(115) and B(119)) xor (A(116) and B(118)) xor (A(117) and B(117)) xor (A(118) and B(116)) xor (A(119) and B(115)) xor (A(120) and B(114)) xor (A(121) and B(113)) xor (A(122) and B(112)) xor (A(123) and B(111)) xor (A(124) and B(110)) xor (A(125) and B(109)) xor (A(126) and B(108)) xor (A(112) and B(127)) xor (A(113) and B(126)) xor (A(114) and B(125)) xor (A(115) and B(124)) xor (A(116) and B(123)) xor (A(117) and B(122)) xor (A(118) and B(121)) xor (A(119) and B(120)) xor (A(120) and B(119)) xor (A(121) and B(118)) xor (A(122) and B(117)) xor (A(123) and B(116)) xor (A(124) and B(115)) xor (A(125) and B(114)) xor (A(126) and B(113)) xor (A(113) and B(127)) xor (A(114) and B(126)) xor (A(115) and B(125)) xor (A(116) and B(124)) xor (A(117) and B(123)) xor (A(118) and B(122)) xor (A(119) and B(121)) xor (A(120) and B(120)) xor (A(121) and B(119)) xor (A(122) and B(118)) xor (A(123) and B(117)) xor (A(124) and B(116)) xor (A(125) and B(115)) xor (A(126) and B(114)) xor (A(114) and B(127)) xor (A(115) and B(126)) xor (A(116) and B(125)) xor (A(117) and B(124)) xor (A(118) and B(123)) xor (A(119) and B(122)) xor (A(120) and B(121)) xor (A(121) and B(120)) xor (A(122) and B(119)) xor (A(123) and B(118)) xor (A(124) and B(117)) xor (A(125) and B(116)) xor (A(126) and B(116));
    C(115) <= (A(0) and B(115)) xor (A(1) and B(114)) xor (A(2) and B(113)) xor (A(3) and B(112)) xor (A(4) and B(111)) xor (A(5) and B(110)) xor (A(6) and B(109)) xor (A(7) and B(108)) xor (A(8) and B(107)) xor (A(9) and B(106)) xor (A(10) and B(105)) xor (A(11) and B(104)) xor (A(12) and B(103)) xor (A(13) and B(102)) xor (A(14) and B(101)) xor (A(15) and B(100)) xor (A(16) and B(99)) xor (A(17) and B(98)) xor (A(18) and B(97)) xor (A(19) and B(96)) xor (A(20) and B(95)) xor (A(21) and B(94)) xor (A(23) and B(93)) xor (A(23) and B(92)) xor (A(24) and B(91)) xor (A(25) and B(90)) xor (A(26) and B(89)) xor (A(27) and B(88)) xor (A(28) and B(87)) xor (A(29) and B(86)) xor (A(30) and B(85)) xor (A(31) and B(84)) xor (A(32) and B(83)) xor (A(33) and B(82)) xor (A(34) and B(81)) xor (A(35) and B(80)) xor (A(36) and B(79)) xor (A(37) and B(78)) xor (A(38) and B(77)) xor (A(39) and B(76)) xor (A(40) and B(75)) xor (A(41) and B(74)) xor (A(42) and B(73)) xor (A(43) and B(72)) xor (A(44) and B(71)) xor (A(45) and B(70)) xor (A(46) and B(69)) xor (A(47) and B(68)) xor (A(48) and B(67)) xor (A(49) and B(66)) xor (A(50) and B(65)) xor (A(51) and B(64)) xor (A(52) and B(63)) xor (A(53) and B(62)) xor (A(54) and B(61)) xor (A(55) and B(60)) xor (A(56) and B(59)) xor (A(57) and B(58)) xor (A(58) and B(57)) xor (A(59) and B(56)) xor (A(60) and B(55)) xor (A(61) and B(54)) xor (A(62) and B(53)) xor (A(63) and B(52)) xor (A(64) and B(51)) xor (A(65) and B(50)) xor (A(66) and B(49)) xor (A(67) and B(48)) xor (A(68) and B(47)) xor (A(69) and B(46)) xor (A(70) and B(45)) xor (A(71) and B(44)) xor (A(72) and B(43)) xor (A(73) and B(42)) xor (A(74) and B(41)) xor (A(75) and B(40)) xor (A(76) and B(39)) xor (A(77) and B(38)) xor (A(78) and B(37)) xor (A(79) and B(36)) xor (A(80) and B(35)) xor (A(81) and B(34)) xor (A(82) and B(33)) xor (A(83) and B(32)) xor (A(84) and B(31)) xor (A(85) and B(30)) xor (A(86) and B(29)) xor (A(87) and B(28)) xor (A(88) and B(27)) xor (A(89) and B(26)) xor (A(90) and B(25)) xor (A(91) and B(24)) xor (A(92) and B(23)) xor (A(93) and B(23)) xor (A(94) and B(21)) xor (A(95) and B(20)) xor (A(96) and B(19)) xor (A(97) and B(18)) xor (A(98) and B(17)) xor (A(99) and B(16)) xor (A(100) and B(15)) xor (A(101) and B(14)) xor (A(102) and B(13)) xor (A(103) and B(12)) xor (A(104) and B(11)) xor (A(105) and B(10)) xor (A(106) and B(9)) xor (A(107) and B(8)) xor (A(108) and B(7)) xor (A(109) and B(6)) xor (A(110) and B(5)) xor (A(111) and B(4)) xor (A(112) and B(3)) xor (A(113) and B(2)) xor (A(114) and B(1)) xor (A(115) and B(0)) xor (A(108) and B(127)) xor (A(109) and B(126)) xor (A(110) and B(125)) xor (A(111) and B(124)) xor (A(112) and B(123)) xor (A(113) and B(122)) xor (A(114) and B(121)) xor (A(115) and B(120)) xor (A(116) and B(119)) xor (A(117) and B(118)) xor (A(118) and B(117)) xor (A(119) and B(116)) xor (A(120) and B(115)) xor (A(121) and B(114)) xor (A(122) and B(113)) xor (A(123) and B(112)) xor (A(124) and B(111)) xor (A(125) and B(110)) xor (A(126) and B(109)) xor (A(113) and B(127)) xor (A(114) and B(126)) xor (A(115) and B(125)) xor (A(116) and B(124)) xor (A(117) and B(123)) xor (A(118) and B(122)) xor (A(119) and B(121)) xor (A(120) and B(120)) xor (A(121) and B(119)) xor (A(122) and B(118)) xor (A(123) and B(117)) xor (A(124) and B(116)) xor (A(125) and B(115)) xor (A(126) and B(114)) xor (A(114) and B(127)) xor (A(115) and B(126)) xor (A(116) and B(125)) xor (A(117) and B(124)) xor (A(118) and B(123)) xor (A(119) and B(122)) xor (A(120) and B(121)) xor (A(121) and B(120)) xor (A(122) and B(119)) xor (A(123) and B(118)) xor (A(124) and B(117)) xor (A(125) and B(116)) xor (A(126) and B(115)) xor (A(115) and B(127)) xor (A(116) and B(126)) xor (A(117) and B(125)) xor (A(118) and B(124)) xor (A(119) and B(123)) xor (A(120) and B(122)) xor (A(121) and B(121)) xor (A(122) and B(120)) xor (A(123) and B(119)) xor (A(124) and B(118)) xor (A(125) and B(117)) xor (A(126) and B(117));
    C(116) <= (A(0) and B(116)) xor (A(1) and B(115)) xor (A(2) and B(114)) xor (A(3) and B(113)) xor (A(4) and B(112)) xor (A(5) and B(111)) xor (A(6) and B(110)) xor (A(7) and B(109)) xor (A(8) and B(108)) xor (A(9) and B(107)) xor (A(10) and B(106)) xor (A(11) and B(105)) xor (A(12) and B(104)) xor (A(13) and B(103)) xor (A(14) and B(102)) xor (A(15) and B(101)) xor (A(16) and B(100)) xor (A(17) and B(99)) xor (A(18) and B(98)) xor (A(19) and B(97)) xor (A(20) and B(96)) xor (A(21) and B(95)) xor (A(23) and B(94)) xor (A(23) and B(93)) xor (A(24) and B(92)) xor (A(25) and B(91)) xor (A(26) and B(90)) xor (A(27) and B(89)) xor (A(28) and B(88)) xor (A(29) and B(87)) xor (A(30) and B(86)) xor (A(31) and B(85)) xor (A(32) and B(84)) xor (A(33) and B(83)) xor (A(34) and B(82)) xor (A(35) and B(81)) xor (A(36) and B(80)) xor (A(37) and B(79)) xor (A(38) and B(78)) xor (A(39) and B(77)) xor (A(40) and B(76)) xor (A(41) and B(75)) xor (A(42) and B(74)) xor (A(43) and B(73)) xor (A(44) and B(72)) xor (A(45) and B(71)) xor (A(46) and B(70)) xor (A(47) and B(69)) xor (A(48) and B(68)) xor (A(49) and B(67)) xor (A(50) and B(66)) xor (A(51) and B(65)) xor (A(52) and B(64)) xor (A(53) and B(63)) xor (A(54) and B(62)) xor (A(55) and B(61)) xor (A(56) and B(60)) xor (A(57) and B(59)) xor (A(58) and B(58)) xor (A(59) and B(57)) xor (A(60) and B(56)) xor (A(61) and B(55)) xor (A(62) and B(54)) xor (A(63) and B(53)) xor (A(64) and B(52)) xor (A(65) and B(51)) xor (A(66) and B(50)) xor (A(67) and B(49)) xor (A(68) and B(48)) xor (A(69) and B(47)) xor (A(70) and B(46)) xor (A(71) and B(45)) xor (A(72) and B(44)) xor (A(73) and B(43)) xor (A(74) and B(42)) xor (A(75) and B(41)) xor (A(76) and B(40)) xor (A(77) and B(39)) xor (A(78) and B(38)) xor (A(79) and B(37)) xor (A(80) and B(36)) xor (A(81) and B(35)) xor (A(82) and B(34)) xor (A(83) and B(33)) xor (A(84) and B(32)) xor (A(85) and B(31)) xor (A(86) and B(30)) xor (A(87) and B(29)) xor (A(88) and B(28)) xor (A(89) and B(27)) xor (A(90) and B(26)) xor (A(91) and B(25)) xor (A(92) and B(24)) xor (A(93) and B(23)) xor (A(94) and B(23)) xor (A(95) and B(21)) xor (A(96) and B(20)) xor (A(97) and B(19)) xor (A(98) and B(18)) xor (A(99) and B(17)) xor (A(100) and B(16)) xor (A(101) and B(15)) xor (A(102) and B(14)) xor (A(103) and B(13)) xor (A(104) and B(12)) xor (A(105) and B(11)) xor (A(106) and B(10)) xor (A(107) and B(9)) xor (A(108) and B(8)) xor (A(109) and B(7)) xor (A(110) and B(6)) xor (A(111) and B(5)) xor (A(112) and B(4)) xor (A(113) and B(3)) xor (A(114) and B(2)) xor (A(115) and B(1)) xor (A(116) and B(0)) xor (A(109) and B(127)) xor (A(110) and B(126)) xor (A(111) and B(125)) xor (A(112) and B(124)) xor (A(113) and B(123)) xor (A(114) and B(122)) xor (A(115) and B(121)) xor (A(116) and B(120)) xor (A(117) and B(119)) xor (A(118) and B(118)) xor (A(119) and B(117)) xor (A(120) and B(116)) xor (A(121) and B(115)) xor (A(122) and B(114)) xor (A(123) and B(113)) xor (A(124) and B(112)) xor (A(125) and B(111)) xor (A(126) and B(110)) xor (A(114) and B(127)) xor (A(115) and B(126)) xor (A(116) and B(125)) xor (A(117) and B(124)) xor (A(118) and B(123)) xor (A(119) and B(122)) xor (A(120) and B(121)) xor (A(121) and B(120)) xor (A(122) and B(119)) xor (A(123) and B(118)) xor (A(124) and B(117)) xor (A(125) and B(116)) xor (A(126) and B(115)) xor (A(115) and B(127)) xor (A(116) and B(126)) xor (A(117) and B(125)) xor (A(118) and B(124)) xor (A(119) and B(123)) xor (A(120) and B(122)) xor (A(121) and B(121)) xor (A(122) and B(120)) xor (A(123) and B(119)) xor (A(124) and B(118)) xor (A(125) and B(117)) xor (A(126) and B(116)) xor (A(116) and B(127)) xor (A(117) and B(126)) xor (A(118) and B(125)) xor (A(119) and B(124)) xor (A(120) and B(123)) xor (A(121) and B(122)) xor (A(122) and B(121)) xor (A(123) and B(120)) xor (A(124) and B(119)) xor (A(125) and B(118)) xor (A(126) and B(118));
    C(117) <= (A(0) and B(117)) xor (A(1) and B(116)) xor (A(2) and B(115)) xor (A(3) and B(114)) xor (A(4) and B(113)) xor (A(5) and B(112)) xor (A(6) and B(111)) xor (A(7) and B(110)) xor (A(8) and B(109)) xor (A(9) and B(108)) xor (A(10) and B(107)) xor (A(11) and B(106)) xor (A(12) and B(105)) xor (A(13) and B(104)) xor (A(14) and B(103)) xor (A(15) and B(102)) xor (A(16) and B(101)) xor (A(17) and B(100)) xor (A(18) and B(99)) xor (A(19) and B(98)) xor (A(20) and B(97)) xor (A(21) and B(96)) xor (A(23) and B(95)) xor (A(23) and B(94)) xor (A(24) and B(93)) xor (A(25) and B(92)) xor (A(26) and B(91)) xor (A(27) and B(90)) xor (A(28) and B(89)) xor (A(29) and B(88)) xor (A(30) and B(87)) xor (A(31) and B(86)) xor (A(32) and B(85)) xor (A(33) and B(84)) xor (A(34) and B(83)) xor (A(35) and B(82)) xor (A(36) and B(81)) xor (A(37) and B(80)) xor (A(38) and B(79)) xor (A(39) and B(78)) xor (A(40) and B(77)) xor (A(41) and B(76)) xor (A(42) and B(75)) xor (A(43) and B(74)) xor (A(44) and B(73)) xor (A(45) and B(72)) xor (A(46) and B(71)) xor (A(47) and B(70)) xor (A(48) and B(69)) xor (A(49) and B(68)) xor (A(50) and B(67)) xor (A(51) and B(66)) xor (A(52) and B(65)) xor (A(53) and B(64)) xor (A(54) and B(63)) xor (A(55) and B(62)) xor (A(56) and B(61)) xor (A(57) and B(60)) xor (A(58) and B(59)) xor (A(59) and B(58)) xor (A(60) and B(57)) xor (A(61) and B(56)) xor (A(62) and B(55)) xor (A(63) and B(54)) xor (A(64) and B(53)) xor (A(65) and B(52)) xor (A(66) and B(51)) xor (A(67) and B(50)) xor (A(68) and B(49)) xor (A(69) and B(48)) xor (A(70) and B(47)) xor (A(71) and B(46)) xor (A(72) and B(45)) xor (A(73) and B(44)) xor (A(74) and B(43)) xor (A(75) and B(42)) xor (A(76) and B(41)) xor (A(77) and B(40)) xor (A(78) and B(39)) xor (A(79) and B(38)) xor (A(80) and B(37)) xor (A(81) and B(36)) xor (A(82) and B(35)) xor (A(83) and B(34)) xor (A(84) and B(33)) xor (A(85) and B(32)) xor (A(86) and B(31)) xor (A(87) and B(30)) xor (A(88) and B(29)) xor (A(89) and B(28)) xor (A(90) and B(27)) xor (A(91) and B(26)) xor (A(92) and B(25)) xor (A(93) and B(24)) xor (A(94) and B(23)) xor (A(95) and B(23)) xor (A(96) and B(21)) xor (A(97) and B(20)) xor (A(98) and B(19)) xor (A(99) and B(18)) xor (A(100) and B(17)) xor (A(101) and B(16)) xor (A(102) and B(15)) xor (A(103) and B(14)) xor (A(104) and B(13)) xor (A(105) and B(12)) xor (A(106) and B(11)) xor (A(107) and B(10)) xor (A(108) and B(9)) xor (A(109) and B(8)) xor (A(110) and B(7)) xor (A(111) and B(6)) xor (A(112) and B(5)) xor (A(113) and B(4)) xor (A(114) and B(3)) xor (A(115) and B(2)) xor (A(116) and B(1)) xor (A(117) and B(0)) xor (A(110) and B(127)) xor (A(111) and B(126)) xor (A(112) and B(125)) xor (A(113) and B(124)) xor (A(114) and B(123)) xor (A(115) and B(122)) xor (A(116) and B(121)) xor (A(117) and B(120)) xor (A(118) and B(119)) xor (A(119) and B(118)) xor (A(120) and B(117)) xor (A(121) and B(116)) xor (A(122) and B(115)) xor (A(123) and B(114)) xor (A(124) and B(113)) xor (A(125) and B(112)) xor (A(126) and B(111)) xor (A(115) and B(127)) xor (A(116) and B(126)) xor (A(117) and B(125)) xor (A(118) and B(124)) xor (A(119) and B(123)) xor (A(120) and B(122)) xor (A(121) and B(121)) xor (A(122) and B(120)) xor (A(123) and B(119)) xor (A(124) and B(118)) xor (A(125) and B(117)) xor (A(126) and B(116)) xor (A(116) and B(127)) xor (A(117) and B(126)) xor (A(118) and B(125)) xor (A(119) and B(124)) xor (A(120) and B(123)) xor (A(121) and B(122)) xor (A(122) and B(121)) xor (A(123) and B(120)) xor (A(124) and B(119)) xor (A(125) and B(118)) xor (A(126) and B(117)) xor (A(117) and B(127)) xor (A(118) and B(126)) xor (A(119) and B(125)) xor (A(120) and B(124)) xor (A(121) and B(123)) xor (A(122) and B(122)) xor (A(123) and B(121)) xor (A(124) and B(120)) xor (A(125) and B(119)) xor (A(126) and B(119));
    C(118) <= (A(0) and B(118)) xor (A(1) and B(117)) xor (A(2) and B(116)) xor (A(3) and B(115)) xor (A(4) and B(114)) xor (A(5) and B(113)) xor (A(6) and B(112)) xor (A(7) and B(111)) xor (A(8) and B(110)) xor (A(9) and B(109)) xor (A(10) and B(108)) xor (A(11) and B(107)) xor (A(12) and B(106)) xor (A(13) and B(105)) xor (A(14) and B(104)) xor (A(15) and B(103)) xor (A(16) and B(102)) xor (A(17) and B(101)) xor (A(18) and B(100)) xor (A(19) and B(99)) xor (A(20) and B(98)) xor (A(21) and B(97)) xor (A(23) and B(96)) xor (A(23) and B(95)) xor (A(24) and B(94)) xor (A(25) and B(93)) xor (A(26) and B(92)) xor (A(27) and B(91)) xor (A(28) and B(90)) xor (A(29) and B(89)) xor (A(30) and B(88)) xor (A(31) and B(87)) xor (A(32) and B(86)) xor (A(33) and B(85)) xor (A(34) and B(84)) xor (A(35) and B(83)) xor (A(36) and B(82)) xor (A(37) and B(81)) xor (A(38) and B(80)) xor (A(39) and B(79)) xor (A(40) and B(78)) xor (A(41) and B(77)) xor (A(42) and B(76)) xor (A(43) and B(75)) xor (A(44) and B(74)) xor (A(45) and B(73)) xor (A(46) and B(72)) xor (A(47) and B(71)) xor (A(48) and B(70)) xor (A(49) and B(69)) xor (A(50) and B(68)) xor (A(51) and B(67)) xor (A(52) and B(66)) xor (A(53) and B(65)) xor (A(54) and B(64)) xor (A(55) and B(63)) xor (A(56) and B(62)) xor (A(57) and B(61)) xor (A(58) and B(60)) xor (A(59) and B(59)) xor (A(60) and B(58)) xor (A(61) and B(57)) xor (A(62) and B(56)) xor (A(63) and B(55)) xor (A(64) and B(54)) xor (A(65) and B(53)) xor (A(66) and B(52)) xor (A(67) and B(51)) xor (A(68) and B(50)) xor (A(69) and B(49)) xor (A(70) and B(48)) xor (A(71) and B(47)) xor (A(72) and B(46)) xor (A(73) and B(45)) xor (A(74) and B(44)) xor (A(75) and B(43)) xor (A(76) and B(42)) xor (A(77) and B(41)) xor (A(78) and B(40)) xor (A(79) and B(39)) xor (A(80) and B(38)) xor (A(81) and B(37)) xor (A(82) and B(36)) xor (A(83) and B(35)) xor (A(84) and B(34)) xor (A(85) and B(33)) xor (A(86) and B(32)) xor (A(87) and B(31)) xor (A(88) and B(30)) xor (A(89) and B(29)) xor (A(90) and B(28)) xor (A(91) and B(27)) xor (A(92) and B(26)) xor (A(93) and B(25)) xor (A(94) and B(24)) xor (A(95) and B(23)) xor (A(96) and B(23)) xor (A(97) and B(21)) xor (A(98) and B(20)) xor (A(99) and B(19)) xor (A(100) and B(18)) xor (A(101) and B(17)) xor (A(102) and B(16)) xor (A(103) and B(15)) xor (A(104) and B(14)) xor (A(105) and B(13)) xor (A(106) and B(12)) xor (A(107) and B(11)) xor (A(108) and B(10)) xor (A(109) and B(9)) xor (A(110) and B(8)) xor (A(111) and B(7)) xor (A(112) and B(6)) xor (A(113) and B(5)) xor (A(114) and B(4)) xor (A(115) and B(3)) xor (A(116) and B(2)) xor (A(117) and B(1)) xor (A(118) and B(0)) xor (A(111) and B(127)) xor (A(112) and B(126)) xor (A(113) and B(125)) xor (A(114) and B(124)) xor (A(115) and B(123)) xor (A(116) and B(122)) xor (A(117) and B(121)) xor (A(118) and B(120)) xor (A(119) and B(119)) xor (A(120) and B(118)) xor (A(121) and B(117)) xor (A(122) and B(116)) xor (A(123) and B(115)) xor (A(124) and B(114)) xor (A(125) and B(113)) xor (A(126) and B(112)) xor (A(116) and B(127)) xor (A(117) and B(126)) xor (A(118) and B(125)) xor (A(119) and B(124)) xor (A(120) and B(123)) xor (A(121) and B(122)) xor (A(122) and B(121)) xor (A(123) and B(120)) xor (A(124) and B(119)) xor (A(125) and B(118)) xor (A(126) and B(117)) xor (A(117) and B(127)) xor (A(118) and B(126)) xor (A(119) and B(125)) xor (A(120) and B(124)) xor (A(121) and B(123)) xor (A(122) and B(122)) xor (A(123) and B(121)) xor (A(124) and B(120)) xor (A(125) and B(119)) xor (A(126) and B(118)) xor (A(118) and B(127)) xor (A(119) and B(126)) xor (A(120) and B(125)) xor (A(121) and B(124)) xor (A(122) and B(123)) xor (A(123) and B(122)) xor (A(124) and B(121)) xor (A(125) and B(120)) xor (A(126) and B(120));
    C(119) <= (A(0) and B(119)) xor (A(1) and B(118)) xor (A(2) and B(117)) xor (A(3) and B(116)) xor (A(4) and B(115)) xor (A(5) and B(114)) xor (A(6) and B(113)) xor (A(7) and B(112)) xor (A(8) and B(111)) xor (A(9) and B(110)) xor (A(10) and B(109)) xor (A(11) and B(108)) xor (A(12) and B(107)) xor (A(13) and B(106)) xor (A(14) and B(105)) xor (A(15) and B(104)) xor (A(16) and B(103)) xor (A(17) and B(102)) xor (A(18) and B(101)) xor (A(19) and B(100)) xor (A(20) and B(99)) xor (A(21) and B(98)) xor (A(23) and B(97)) xor (A(23) and B(96)) xor (A(24) and B(95)) xor (A(25) and B(94)) xor (A(26) and B(93)) xor (A(27) and B(92)) xor (A(28) and B(91)) xor (A(29) and B(90)) xor (A(30) and B(89)) xor (A(31) and B(88)) xor (A(32) and B(87)) xor (A(33) and B(86)) xor (A(34) and B(85)) xor (A(35) and B(84)) xor (A(36) and B(83)) xor (A(37) and B(82)) xor (A(38) and B(81)) xor (A(39) and B(80)) xor (A(40) and B(79)) xor (A(41) and B(78)) xor (A(42) and B(77)) xor (A(43) and B(76)) xor (A(44) and B(75)) xor (A(45) and B(74)) xor (A(46) and B(73)) xor (A(47) and B(72)) xor (A(48) and B(71)) xor (A(49) and B(70)) xor (A(50) and B(69)) xor (A(51) and B(68)) xor (A(52) and B(67)) xor (A(53) and B(66)) xor (A(54) and B(65)) xor (A(55) and B(64)) xor (A(56) and B(63)) xor (A(57) and B(62)) xor (A(58) and B(61)) xor (A(59) and B(60)) xor (A(60) and B(59)) xor (A(61) and B(58)) xor (A(62) and B(57)) xor (A(63) and B(56)) xor (A(64) and B(55)) xor (A(65) and B(54)) xor (A(66) and B(53)) xor (A(67) and B(52)) xor (A(68) and B(51)) xor (A(69) and B(50)) xor (A(70) and B(49)) xor (A(71) and B(48)) xor (A(72) and B(47)) xor (A(73) and B(46)) xor (A(74) and B(45)) xor (A(75) and B(44)) xor (A(76) and B(43)) xor (A(77) and B(42)) xor (A(78) and B(41)) xor (A(79) and B(40)) xor (A(80) and B(39)) xor (A(81) and B(38)) xor (A(82) and B(37)) xor (A(83) and B(36)) xor (A(84) and B(35)) xor (A(85) and B(34)) xor (A(86) and B(33)) xor (A(87) and B(32)) xor (A(88) and B(31)) xor (A(89) and B(30)) xor (A(90) and B(29)) xor (A(91) and B(28)) xor (A(92) and B(27)) xor (A(93) and B(26)) xor (A(94) and B(25)) xor (A(95) and B(24)) xor (A(96) and B(23)) xor (A(97) and B(23)) xor (A(98) and B(21)) xor (A(99) and B(20)) xor (A(100) and B(19)) xor (A(101) and B(18)) xor (A(102) and B(17)) xor (A(103) and B(16)) xor (A(104) and B(15)) xor (A(105) and B(14)) xor (A(106) and B(13)) xor (A(107) and B(12)) xor (A(108) and B(11)) xor (A(109) and B(10)) xor (A(110) and B(9)) xor (A(111) and B(8)) xor (A(112) and B(7)) xor (A(113) and B(6)) xor (A(114) and B(5)) xor (A(115) and B(4)) xor (A(116) and B(3)) xor (A(117) and B(2)) xor (A(118) and B(1)) xor (A(119) and B(0)) xor (A(112) and B(127)) xor (A(113) and B(126)) xor (A(114) and B(125)) xor (A(115) and B(124)) xor (A(116) and B(123)) xor (A(117) and B(122)) xor (A(118) and B(121)) xor (A(119) and B(120)) xor (A(120) and B(119)) xor (A(121) and B(118)) xor (A(122) and B(117)) xor (A(123) and B(116)) xor (A(124) and B(115)) xor (A(125) and B(114)) xor (A(126) and B(113)) xor (A(117) and B(127)) xor (A(118) and B(126)) xor (A(119) and B(125)) xor (A(120) and B(124)) xor (A(121) and B(123)) xor (A(122) and B(122)) xor (A(123) and B(121)) xor (A(124) and B(120)) xor (A(125) and B(119)) xor (A(126) and B(118)) xor (A(118) and B(127)) xor (A(119) and B(126)) xor (A(120) and B(125)) xor (A(121) and B(124)) xor (A(122) and B(123)) xor (A(123) and B(122)) xor (A(124) and B(121)) xor (A(125) and B(120)) xor (A(126) and B(119)) xor (A(119) and B(127)) xor (A(120) and B(126)) xor (A(121) and B(125)) xor (A(122) and B(124)) xor (A(123) and B(123)) xor (A(124) and B(122)) xor (A(125) and B(121)) xor (A(126) and B(121));
    C(120) <= (A(0) and B(120)) xor (A(1) and B(119)) xor (A(2) and B(118)) xor (A(3) and B(117)) xor (A(4) and B(116)) xor (A(5) and B(115)) xor (A(6) and B(114)) xor (A(7) and B(113)) xor (A(8) and B(112)) xor (A(9) and B(111)) xor (A(10) and B(110)) xor (A(11) and B(109)) xor (A(12) and B(108)) xor (A(13) and B(107)) xor (A(14) and B(106)) xor (A(15) and B(105)) xor (A(16) and B(104)) xor (A(17) and B(103)) xor (A(18) and B(102)) xor (A(19) and B(101)) xor (A(20) and B(100)) xor (A(21) and B(99)) xor (A(23) and B(98)) xor (A(23) and B(97)) xor (A(24) and B(96)) xor (A(25) and B(95)) xor (A(26) and B(94)) xor (A(27) and B(93)) xor (A(28) and B(92)) xor (A(29) and B(91)) xor (A(30) and B(90)) xor (A(31) and B(89)) xor (A(32) and B(88)) xor (A(33) and B(87)) xor (A(34) and B(86)) xor (A(35) and B(85)) xor (A(36) and B(84)) xor (A(37) and B(83)) xor (A(38) and B(82)) xor (A(39) and B(81)) xor (A(40) and B(80)) xor (A(41) and B(79)) xor (A(42) and B(78)) xor (A(43) and B(77)) xor (A(44) and B(76)) xor (A(45) and B(75)) xor (A(46) and B(74)) xor (A(47) and B(73)) xor (A(48) and B(72)) xor (A(49) and B(71)) xor (A(50) and B(70)) xor (A(51) and B(69)) xor (A(52) and B(68)) xor (A(53) and B(67)) xor (A(54) and B(66)) xor (A(55) and B(65)) xor (A(56) and B(64)) xor (A(57) and B(63)) xor (A(58) and B(62)) xor (A(59) and B(61)) xor (A(60) and B(60)) xor (A(61) and B(59)) xor (A(62) and B(58)) xor (A(63) and B(57)) xor (A(64) and B(56)) xor (A(65) and B(55)) xor (A(66) and B(54)) xor (A(67) and B(53)) xor (A(68) and B(52)) xor (A(69) and B(51)) xor (A(70) and B(50)) xor (A(71) and B(49)) xor (A(72) and B(48)) xor (A(73) and B(47)) xor (A(74) and B(46)) xor (A(75) and B(45)) xor (A(76) and B(44)) xor (A(77) and B(43)) xor (A(78) and B(42)) xor (A(79) and B(41)) xor (A(80) and B(40)) xor (A(81) and B(39)) xor (A(82) and B(38)) xor (A(83) and B(37)) xor (A(84) and B(36)) xor (A(85) and B(35)) xor (A(86) and B(34)) xor (A(87) and B(33)) xor (A(88) and B(32)) xor (A(89) and B(31)) xor (A(90) and B(30)) xor (A(91) and B(29)) xor (A(92) and B(28)) xor (A(93) and B(27)) xor (A(94) and B(26)) xor (A(95) and B(25)) xor (A(96) and B(24)) xor (A(97) and B(23)) xor (A(98) and B(23)) xor (A(99) and B(21)) xor (A(100) and B(20)) xor (A(101) and B(19)) xor (A(102) and B(18)) xor (A(103) and B(17)) xor (A(104) and B(16)) xor (A(105) and B(15)) xor (A(106) and B(14)) xor (A(107) and B(13)) xor (A(108) and B(12)) xor (A(109) and B(11)) xor (A(110) and B(10)) xor (A(111) and B(9)) xor (A(112) and B(8)) xor (A(113) and B(7)) xor (A(114) and B(6)) xor (A(115) and B(5)) xor (A(116) and B(4)) xor (A(117) and B(3)) xor (A(118) and B(2)) xor (A(119) and B(1)) xor (A(120) and B(0)) xor (A(113) and B(127)) xor (A(114) and B(126)) xor (A(115) and B(125)) xor (A(116) and B(124)) xor (A(117) and B(123)) xor (A(118) and B(122)) xor (A(119) and B(121)) xor (A(120) and B(120)) xor (A(121) and B(119)) xor (A(122) and B(118)) xor (A(123) and B(117)) xor (A(124) and B(116)) xor (A(125) and B(115)) xor (A(126) and B(114)) xor (A(118) and B(127)) xor (A(119) and B(126)) xor (A(120) and B(125)) xor (A(121) and B(124)) xor (A(122) and B(123)) xor (A(123) and B(122)) xor (A(124) and B(121)) xor (A(125) and B(120)) xor (A(126) and B(119)) xor (A(119) and B(127)) xor (A(120) and B(126)) xor (A(121) and B(125)) xor (A(122) and B(124)) xor (A(123) and B(123)) xor (A(124) and B(122)) xor (A(125) and B(121)) xor (A(126) and B(120)) xor (A(120) and B(127)) xor (A(121) and B(126)) xor (A(122) and B(125)) xor (A(123) and B(124)) xor (A(124) and B(123)) xor (A(125) and B(122)) xor (A(126) and B(122));
    C(121) <= (A(0) and B(121)) xor (A(1) and B(120)) xor (A(2) and B(119)) xor (A(3) and B(118)) xor (A(4) and B(117)) xor (A(5) and B(116)) xor (A(6) and B(115)) xor (A(7) and B(114)) xor (A(8) and B(113)) xor (A(9) and B(112)) xor (A(10) and B(111)) xor (A(11) and B(110)) xor (A(12) and B(109)) xor (A(13) and B(108)) xor (A(14) and B(107)) xor (A(15) and B(106)) xor (A(16) and B(105)) xor (A(17) and B(104)) xor (A(18) and B(103)) xor (A(19) and B(102)) xor (A(20) and B(101)) xor (A(21) and B(100)) xor (A(23) and B(99)) xor (A(23) and B(98)) xor (A(24) and B(97)) xor (A(25) and B(96)) xor (A(26) and B(95)) xor (A(27) and B(94)) xor (A(28) and B(93)) xor (A(29) and B(92)) xor (A(30) and B(91)) xor (A(31) and B(90)) xor (A(32) and B(89)) xor (A(33) and B(88)) xor (A(34) and B(87)) xor (A(35) and B(86)) xor (A(36) and B(85)) xor (A(37) and B(84)) xor (A(38) and B(83)) xor (A(39) and B(82)) xor (A(40) and B(81)) xor (A(41) and B(80)) xor (A(42) and B(79)) xor (A(43) and B(78)) xor (A(44) and B(77)) xor (A(45) and B(76)) xor (A(46) and B(75)) xor (A(47) and B(74)) xor (A(48) and B(73)) xor (A(49) and B(72)) xor (A(50) and B(71)) xor (A(51) and B(70)) xor (A(52) and B(69)) xor (A(53) and B(68)) xor (A(54) and B(67)) xor (A(55) and B(66)) xor (A(56) and B(65)) xor (A(57) and B(64)) xor (A(58) and B(63)) xor (A(59) and B(62)) xor (A(60) and B(61)) xor (A(61) and B(60)) xor (A(62) and B(59)) xor (A(63) and B(58)) xor (A(64) and B(57)) xor (A(65) and B(56)) xor (A(66) and B(55)) xor (A(67) and B(54)) xor (A(68) and B(53)) xor (A(69) and B(52)) xor (A(70) and B(51)) xor (A(71) and B(50)) xor (A(72) and B(49)) xor (A(73) and B(48)) xor (A(74) and B(47)) xor (A(75) and B(46)) xor (A(76) and B(45)) xor (A(77) and B(44)) xor (A(78) and B(43)) xor (A(79) and B(42)) xor (A(80) and B(41)) xor (A(81) and B(40)) xor (A(82) and B(39)) xor (A(83) and B(38)) xor (A(84) and B(37)) xor (A(85) and B(36)) xor (A(86) and B(35)) xor (A(87) and B(34)) xor (A(88) and B(33)) xor (A(89) and B(32)) xor (A(90) and B(31)) xor (A(91) and B(30)) xor (A(92) and B(29)) xor (A(93) and B(28)) xor (A(94) and B(27)) xor (A(95) and B(26)) xor (A(96) and B(25)) xor (A(97) and B(24)) xor (A(98) and B(23)) xor (A(99) and B(23)) xor (A(100) and B(21)) xor (A(101) and B(20)) xor (A(102) and B(19)) xor (A(103) and B(18)) xor (A(104) and B(17)) xor (A(105) and B(16)) xor (A(106) and B(15)) xor (A(107) and B(14)) xor (A(108) and B(13)) xor (A(109) and B(12)) xor (A(110) and B(11)) xor (A(111) and B(10)) xor (A(112) and B(9)) xor (A(113) and B(8)) xor (A(114) and B(7)) xor (A(115) and B(6)) xor (A(116) and B(5)) xor (A(117) and B(4)) xor (A(118) and B(3)) xor (A(119) and B(2)) xor (A(120) and B(1)) xor (A(121) and B(0)) xor (A(114) and B(127)) xor (A(115) and B(126)) xor (A(116) and B(125)) xor (A(117) and B(124)) xor (A(118) and B(123)) xor (A(119) and B(122)) xor (A(120) and B(121)) xor (A(121) and B(120)) xor (A(122) and B(119)) xor (A(123) and B(118)) xor (A(124) and B(117)) xor (A(125) and B(116)) xor (A(126) and B(115)) xor (A(119) and B(127)) xor (A(120) and B(126)) xor (A(121) and B(125)) xor (A(122) and B(124)) xor (A(123) and B(123)) xor (A(124) and B(122)) xor (A(125) and B(121)) xor (A(126) and B(120)) xor (A(120) and B(127)) xor (A(121) and B(126)) xor (A(122) and B(125)) xor (A(123) and B(124)) xor (A(124) and B(123)) xor (A(125) and B(122)) xor (A(126) and B(121)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(123));
    C(122) <= (A(0) and B(122)) xor (A(1) and B(121)) xor (A(2) and B(120)) xor (A(3) and B(119)) xor (A(4) and B(118)) xor (A(5) and B(117)) xor (A(6) and B(116)) xor (A(7) and B(115)) xor (A(8) and B(114)) xor (A(9) and B(113)) xor (A(10) and B(112)) xor (A(11) and B(111)) xor (A(12) and B(110)) xor (A(13) and B(109)) xor (A(14) and B(108)) xor (A(15) and B(107)) xor (A(16) and B(106)) xor (A(17) and B(105)) xor (A(18) and B(104)) xor (A(19) and B(103)) xor (A(20) and B(102)) xor (A(21) and B(101)) xor (A(23) and B(100)) xor (A(23) and B(99)) xor (A(24) and B(98)) xor (A(25) and B(97)) xor (A(26) and B(96)) xor (A(27) and B(95)) xor (A(28) and B(94)) xor (A(29) and B(93)) xor (A(30) and B(92)) xor (A(31) and B(91)) xor (A(32) and B(90)) xor (A(33) and B(89)) xor (A(34) and B(88)) xor (A(35) and B(87)) xor (A(36) and B(86)) xor (A(37) and B(85)) xor (A(38) and B(84)) xor (A(39) and B(83)) xor (A(40) and B(82)) xor (A(41) and B(81)) xor (A(42) and B(80)) xor (A(43) and B(79)) xor (A(44) and B(78)) xor (A(45) and B(77)) xor (A(46) and B(76)) xor (A(47) and B(75)) xor (A(48) and B(74)) xor (A(49) and B(73)) xor (A(50) and B(72)) xor (A(51) and B(71)) xor (A(52) and B(70)) xor (A(53) and B(69)) xor (A(54) and B(68)) xor (A(55) and B(67)) xor (A(56) and B(66)) xor (A(57) and B(65)) xor (A(58) and B(64)) xor (A(59) and B(63)) xor (A(60) and B(62)) xor (A(61) and B(61)) xor (A(62) and B(60)) xor (A(63) and B(59)) xor (A(64) and B(58)) xor (A(65) and B(57)) xor (A(66) and B(56)) xor (A(67) and B(55)) xor (A(68) and B(54)) xor (A(69) and B(53)) xor (A(70) and B(52)) xor (A(71) and B(51)) xor (A(72) and B(50)) xor (A(73) and B(49)) xor (A(74) and B(48)) xor (A(75) and B(47)) xor (A(76) and B(46)) xor (A(77) and B(45)) xor (A(78) and B(44)) xor (A(79) and B(43)) xor (A(80) and B(42)) xor (A(81) and B(41)) xor (A(82) and B(40)) xor (A(83) and B(39)) xor (A(84) and B(38)) xor (A(85) and B(37)) xor (A(86) and B(36)) xor (A(87) and B(35)) xor (A(88) and B(34)) xor (A(89) and B(33)) xor (A(90) and B(32)) xor (A(91) and B(31)) xor (A(92) and B(30)) xor (A(93) and B(29)) xor (A(94) and B(28)) xor (A(95) and B(27)) xor (A(96) and B(26)) xor (A(97) and B(25)) xor (A(98) and B(24)) xor (A(99) and B(23)) xor (A(100) and B(23)) xor (A(101) and B(21)) xor (A(102) and B(20)) xor (A(103) and B(19)) xor (A(104) and B(18)) xor (A(105) and B(17)) xor (A(106) and B(16)) xor (A(107) and B(15)) xor (A(108) and B(14)) xor (A(109) and B(13)) xor (A(110) and B(12)) xor (A(111) and B(11)) xor (A(112) and B(10)) xor (A(113) and B(9)) xor (A(114) and B(8)) xor (A(115) and B(7)) xor (A(116) and B(6)) xor (A(117) and B(5)) xor (A(118) and B(4)) xor (A(119) and B(3)) xor (A(120) and B(2)) xor (A(121) and B(1)) xor (A(122) and B(0)) xor (A(115) and B(127)) xor (A(116) and B(126)) xor (A(117) and B(125)) xor (A(118) and B(124)) xor (A(119) and B(123)) xor (A(120) and B(122)) xor (A(121) and B(121)) xor (A(122) and B(120)) xor (A(123) and B(119)) xor (A(124) and B(118)) xor (A(125) and B(117)) xor (A(126) and B(116)) xor (A(120) and B(127)) xor (A(121) and B(126)) xor (A(122) and B(125)) xor (A(123) and B(124)) xor (A(124) and B(123)) xor (A(125) and B(122)) xor (A(126) and B(121)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(122)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(124));
    C(123) <= (A(0) and B(123)) xor (A(1) and B(122)) xor (A(2) and B(121)) xor (A(3) and B(120)) xor (A(4) and B(119)) xor (A(5) and B(118)) xor (A(6) and B(117)) xor (A(7) and B(116)) xor (A(8) and B(115)) xor (A(9) and B(114)) xor (A(10) and B(113)) xor (A(11) and B(112)) xor (A(12) and B(111)) xor (A(13) and B(110)) xor (A(14) and B(109)) xor (A(15) and B(108)) xor (A(16) and B(107)) xor (A(17) and B(106)) xor (A(18) and B(105)) xor (A(19) and B(104)) xor (A(20) and B(103)) xor (A(21) and B(102)) xor (A(23) and B(101)) xor (A(23) and B(100)) xor (A(24) and B(99)) xor (A(25) and B(98)) xor (A(26) and B(97)) xor (A(27) and B(96)) xor (A(28) and B(95)) xor (A(29) and B(94)) xor (A(30) and B(93)) xor (A(31) and B(92)) xor (A(32) and B(91)) xor (A(33) and B(90)) xor (A(34) and B(89)) xor (A(35) and B(88)) xor (A(36) and B(87)) xor (A(37) and B(86)) xor (A(38) and B(85)) xor (A(39) and B(84)) xor (A(40) and B(83)) xor (A(41) and B(82)) xor (A(42) and B(81)) xor (A(43) and B(80)) xor (A(44) and B(79)) xor (A(45) and B(78)) xor (A(46) and B(77)) xor (A(47) and B(76)) xor (A(48) and B(75)) xor (A(49) and B(74)) xor (A(50) and B(73)) xor (A(51) and B(72)) xor (A(52) and B(71)) xor (A(53) and B(70)) xor (A(54) and B(69)) xor (A(55) and B(68)) xor (A(56) and B(67)) xor (A(57) and B(66)) xor (A(58) and B(65)) xor (A(59) and B(64)) xor (A(60) and B(63)) xor (A(61) and B(62)) xor (A(62) and B(61)) xor (A(63) and B(60)) xor (A(64) and B(59)) xor (A(65) and B(58)) xor (A(66) and B(57)) xor (A(67) and B(56)) xor (A(68) and B(55)) xor (A(69) and B(54)) xor (A(70) and B(53)) xor (A(71) and B(52)) xor (A(72) and B(51)) xor (A(73) and B(50)) xor (A(74) and B(49)) xor (A(75) and B(48)) xor (A(76) and B(47)) xor (A(77) and B(46)) xor (A(78) and B(45)) xor (A(79) and B(44)) xor (A(80) and B(43)) xor (A(81) and B(42)) xor (A(82) and B(41)) xor (A(83) and B(40)) xor (A(84) and B(39)) xor (A(85) and B(38)) xor (A(86) and B(37)) xor (A(87) and B(36)) xor (A(88) and B(35)) xor (A(89) and B(34)) xor (A(90) and B(33)) xor (A(91) and B(32)) xor (A(92) and B(31)) xor (A(93) and B(30)) xor (A(94) and B(29)) xor (A(95) and B(28)) xor (A(96) and B(27)) xor (A(97) and B(26)) xor (A(98) and B(25)) xor (A(99) and B(24)) xor (A(100) and B(23)) xor (A(101) and B(23)) xor (A(102) and B(21)) xor (A(103) and B(20)) xor (A(104) and B(19)) xor (A(105) and B(18)) xor (A(106) and B(17)) xor (A(107) and B(16)) xor (A(108) and B(15)) xor (A(109) and B(14)) xor (A(110) and B(13)) xor (A(111) and B(12)) xor (A(112) and B(11)) xor (A(113) and B(10)) xor (A(114) and B(9)) xor (A(115) and B(8)) xor (A(116) and B(7)) xor (A(117) and B(6)) xor (A(118) and B(5)) xor (A(119) and B(4)) xor (A(120) and B(3)) xor (A(121) and B(2)) xor (A(122) and B(1)) xor (A(123) and B(0)) xor (A(116) and B(127)) xor (A(117) and B(126)) xor (A(118) and B(125)) xor (A(119) and B(124)) xor (A(120) and B(123)) xor (A(121) and B(122)) xor (A(122) and B(121)) xor (A(123) and B(120)) xor (A(124) and B(119)) xor (A(125) and B(118)) xor (A(126) and B(117)) xor (A(121) and B(127)) xor (A(122) and B(126)) xor (A(123) and B(125)) xor (A(124) and B(124)) xor (A(125) and B(123)) xor (A(126) and B(122)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(123)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(125));
    C(124) <= (A(0) and B(124)) xor (A(1) and B(123)) xor (A(2) and B(122)) xor (A(3) and B(121)) xor (A(4) and B(120)) xor (A(5) and B(119)) xor (A(6) and B(118)) xor (A(7) and B(117)) xor (A(8) and B(116)) xor (A(9) and B(115)) xor (A(10) and B(114)) xor (A(11) and B(113)) xor (A(12) and B(112)) xor (A(13) and B(111)) xor (A(14) and B(110)) xor (A(15) and B(109)) xor (A(16) and B(108)) xor (A(17) and B(107)) xor (A(18) and B(106)) xor (A(19) and B(105)) xor (A(20) and B(104)) xor (A(21) and B(103)) xor (A(23) and B(102)) xor (A(23) and B(101)) xor (A(24) and B(100)) xor (A(25) and B(99)) xor (A(26) and B(98)) xor (A(27) and B(97)) xor (A(28) and B(96)) xor (A(29) and B(95)) xor (A(30) and B(94)) xor (A(31) and B(93)) xor (A(32) and B(92)) xor (A(33) and B(91)) xor (A(34) and B(90)) xor (A(35) and B(89)) xor (A(36) and B(88)) xor (A(37) and B(87)) xor (A(38) and B(86)) xor (A(39) and B(85)) xor (A(40) and B(84)) xor (A(41) and B(83)) xor (A(42) and B(82)) xor (A(43) and B(81)) xor (A(44) and B(80)) xor (A(45) and B(79)) xor (A(46) and B(78)) xor (A(47) and B(77)) xor (A(48) and B(76)) xor (A(49) and B(75)) xor (A(50) and B(74)) xor (A(51) and B(73)) xor (A(52) and B(72)) xor (A(53) and B(71)) xor (A(54) and B(70)) xor (A(55) and B(69)) xor (A(56) and B(68)) xor (A(57) and B(67)) xor (A(58) and B(66)) xor (A(59) and B(65)) xor (A(60) and B(64)) xor (A(61) and B(63)) xor (A(62) and B(62)) xor (A(63) and B(61)) xor (A(64) and B(60)) xor (A(65) and B(59)) xor (A(66) and B(58)) xor (A(67) and B(57)) xor (A(68) and B(56)) xor (A(69) and B(55)) xor (A(70) and B(54)) xor (A(71) and B(53)) xor (A(72) and B(52)) xor (A(73) and B(51)) xor (A(74) and B(50)) xor (A(75) and B(49)) xor (A(76) and B(48)) xor (A(77) and B(47)) xor (A(78) and B(46)) xor (A(79) and B(45)) xor (A(80) and B(44)) xor (A(81) and B(43)) xor (A(82) and B(42)) xor (A(83) and B(41)) xor (A(84) and B(40)) xor (A(85) and B(39)) xor (A(86) and B(38)) xor (A(87) and B(37)) xor (A(88) and B(36)) xor (A(89) and B(35)) xor (A(90) and B(34)) xor (A(91) and B(33)) xor (A(92) and B(32)) xor (A(93) and B(31)) xor (A(94) and B(30)) xor (A(95) and B(29)) xor (A(96) and B(28)) xor (A(97) and B(27)) xor (A(98) and B(26)) xor (A(99) and B(25)) xor (A(100) and B(24)) xor (A(101) and B(23)) xor (A(102) and B(23)) xor (A(103) and B(21)) xor (A(104) and B(20)) xor (A(105) and B(19)) xor (A(106) and B(18)) xor (A(107) and B(17)) xor (A(108) and B(16)) xor (A(109) and B(15)) xor (A(110) and B(14)) xor (A(111) and B(13)) xor (A(112) and B(12)) xor (A(113) and B(11)) xor (A(114) and B(10)) xor (A(115) and B(9)) xor (A(116) and B(8)) xor (A(117) and B(7)) xor (A(118) and B(6)) xor (A(119) and B(5)) xor (A(120) and B(4)) xor (A(121) and B(3)) xor (A(122) and B(2)) xor (A(123) and B(1)) xor (A(124) and B(0)) xor (A(117) and B(127)) xor (A(118) and B(126)) xor (A(119) and B(125)) xor (A(120) and B(124)) xor (A(121) and B(123)) xor (A(122) and B(122)) xor (A(123) and B(121)) xor (A(124) and B(120)) xor (A(125) and B(119)) xor (A(126) and B(118)) xor (A(122) and B(127)) xor (A(123) and B(126)) xor (A(124) and B(125)) xor (A(125) and B(124)) xor (A(126) and B(123)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(124)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(126));
    C(125) <= (A(0) and B(125)) xor (A(1) and B(124)) xor (A(2) and B(123)) xor (A(3) and B(122)) xor (A(4) and B(121)) xor (A(5) and B(120)) xor (A(6) and B(119)) xor (A(7) and B(118)) xor (A(8) and B(117)) xor (A(9) and B(116)) xor (A(10) and B(115)) xor (A(11) and B(114)) xor (A(12) and B(113)) xor (A(13) and B(112)) xor (A(14) and B(111)) xor (A(15) and B(110)) xor (A(16) and B(109)) xor (A(17) and B(108)) xor (A(18) and B(107)) xor (A(19) and B(106)) xor (A(20) and B(105)) xor (A(21) and B(104)) xor (A(23) and B(103)) xor (A(23) and B(102)) xor (A(24) and B(101)) xor (A(25) and B(100)) xor (A(26) and B(99)) xor (A(27) and B(98)) xor (A(28) and B(97)) xor (A(29) and B(96)) xor (A(30) and B(95)) xor (A(31) and B(94)) xor (A(32) and B(93)) xor (A(33) and B(92)) xor (A(34) and B(91)) xor (A(35) and B(90)) xor (A(36) and B(89)) xor (A(37) and B(88)) xor (A(38) and B(87)) xor (A(39) and B(86)) xor (A(40) and B(85)) xor (A(41) and B(84)) xor (A(42) and B(83)) xor (A(43) and B(82)) xor (A(44) and B(81)) xor (A(45) and B(80)) xor (A(46) and B(79)) xor (A(47) and B(78)) xor (A(48) and B(77)) xor (A(49) and B(76)) xor (A(50) and B(75)) xor (A(51) and B(74)) xor (A(52) and B(73)) xor (A(53) and B(72)) xor (A(54) and B(71)) xor (A(55) and B(70)) xor (A(56) and B(69)) xor (A(57) and B(68)) xor (A(58) and B(67)) xor (A(59) and B(66)) xor (A(60) and B(65)) xor (A(61) and B(64)) xor (A(62) and B(63)) xor (A(63) and B(62)) xor (A(64) and B(61)) xor (A(65) and B(60)) xor (A(66) and B(59)) xor (A(67) and B(58)) xor (A(68) and B(57)) xor (A(69) and B(56)) xor (A(70) and B(55)) xor (A(71) and B(54)) xor (A(72) and B(53)) xor (A(73) and B(52)) xor (A(74) and B(51)) xor (A(75) and B(50)) xor (A(76) and B(49)) xor (A(77) and B(48)) xor (A(78) and B(47)) xor (A(79) and B(46)) xor (A(80) and B(45)) xor (A(81) and B(44)) xor (A(82) and B(43)) xor (A(83) and B(42)) xor (A(84) and B(41)) xor (A(85) and B(40)) xor (A(86) and B(39)) xor (A(87) and B(38)) xor (A(88) and B(37)) xor (A(89) and B(36)) xor (A(90) and B(35)) xor (A(91) and B(34)) xor (A(92) and B(33)) xor (A(93) and B(32)) xor (A(94) and B(31)) xor (A(95) and B(30)) xor (A(96) and B(29)) xor (A(97) and B(28)) xor (A(98) and B(27)) xor (A(99) and B(26)) xor (A(100) and B(25)) xor (A(101) and B(24)) xor (A(102) and B(23)) xor (A(103) and B(23)) xor (A(104) and B(21)) xor (A(105) and B(20)) xor (A(106) and B(19)) xor (A(107) and B(18)) xor (A(108) and B(17)) xor (A(109) and B(16)) xor (A(110) and B(15)) xor (A(111) and B(14)) xor (A(112) and B(13)) xor (A(113) and B(12)) xor (A(114) and B(11)) xor (A(115) and B(10)) xor (A(116) and B(9)) xor (A(117) and B(8)) xor (A(118) and B(7)) xor (A(119) and B(6)) xor (A(120) and B(5)) xor (A(121) and B(4)) xor (A(122) and B(3)) xor (A(123) and B(2)) xor (A(124) and B(1)) xor (A(125) and B(0)) xor (A(118) and B(127)) xor (A(119) and B(126)) xor (A(120) and B(125)) xor (A(121) and B(124)) xor (A(122) and B(123)) xor (A(123) and B(122)) xor (A(124) and B(121)) xor (A(125) and B(120)) xor (A(126) and B(119)) xor (A(123) and B(127)) xor (A(124) and B(126)) xor (A(125) and B(125)) xor (A(126) and B(124)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(125)) xor (A(125) and B(127)) xor (A(126) and B(127));
    C(126) <= (A(0) and B(126)) xor (A(1) and B(125)) xor (A(2) and B(124)) xor (A(3) and B(123)) xor (A(4) and B(122)) xor (A(5) and B(121)) xor (A(6) and B(120)) xor (A(7) and B(119)) xor (A(8) and B(118)) xor (A(9) and B(117)) xor (A(10) and B(116)) xor (A(11) and B(115)) xor (A(12) and B(114)) xor (A(13) and B(113)) xor (A(14) and B(112)) xor (A(15) and B(111)) xor (A(16) and B(110)) xor (A(17) and B(109)) xor (A(18) and B(108)) xor (A(19) and B(107)) xor (A(20) and B(106)) xor (A(21) and B(105)) xor (A(23) and B(104)) xor (A(23) and B(103)) xor (A(24) and B(102)) xor (A(25) and B(101)) xor (A(26) and B(100)) xor (A(27) and B(99)) xor (A(28) and B(98)) xor (A(29) and B(97)) xor (A(30) and B(96)) xor (A(31) and B(95)) xor (A(32) and B(94)) xor (A(33) and B(93)) xor (A(34) and B(92)) xor (A(35) and B(91)) xor (A(36) and B(90)) xor (A(37) and B(89)) xor (A(38) and B(88)) xor (A(39) and B(87)) xor (A(40) and B(86)) xor (A(41) and B(85)) xor (A(42) and B(84)) xor (A(43) and B(83)) xor (A(44) and B(82)) xor (A(45) and B(81)) xor (A(46) and B(80)) xor (A(47) and B(79)) xor (A(48) and B(78)) xor (A(49) and B(77)) xor (A(50) and B(76)) xor (A(51) and B(75)) xor (A(52) and B(74)) xor (A(53) and B(73)) xor (A(54) and B(72)) xor (A(55) and B(71)) xor (A(56) and B(70)) xor (A(57) and B(69)) xor (A(58) and B(68)) xor (A(59) and B(67)) xor (A(60) and B(66)) xor (A(61) and B(65)) xor (A(62) and B(64)) xor (A(63) and B(63)) xor (A(64) and B(62)) xor (A(65) and B(61)) xor (A(66) and B(60)) xor (A(67) and B(59)) xor (A(68) and B(58)) xor (A(69) and B(57)) xor (A(70) and B(56)) xor (A(71) and B(55)) xor (A(72) and B(54)) xor (A(73) and B(53)) xor (A(74) and B(52)) xor (A(75) and B(51)) xor (A(76) and B(50)) xor (A(77) and B(49)) xor (A(78) and B(48)) xor (A(79) and B(47)) xor (A(80) and B(46)) xor (A(81) and B(45)) xor (A(82) and B(44)) xor (A(83) and B(43)) xor (A(84) and B(42)) xor (A(85) and B(41)) xor (A(86) and B(40)) xor (A(87) and B(39)) xor (A(88) and B(38)) xor (A(89) and B(37)) xor (A(90) and B(36)) xor (A(91) and B(35)) xor (A(92) and B(34)) xor (A(93) and B(33)) xor (A(94) and B(32)) xor (A(95) and B(31)) xor (A(96) and B(30)) xor (A(97) and B(29)) xor (A(98) and B(28)) xor (A(99) and B(27)) xor (A(100) and B(26)) xor (A(101) and B(25)) xor (A(102) and B(24)) xor (A(103) and B(23)) xor (A(104) and B(23)) xor (A(105) and B(21)) xor (A(106) and B(20)) xor (A(107) and B(19)) xor (A(108) and B(18)) xor (A(109) and B(17)) xor (A(110) and B(16)) xor (A(111) and B(15)) xor (A(112) and B(14)) xor (A(113) and B(13)) xor (A(114) and B(12)) xor (A(115) and B(11)) xor (A(116) and B(10)) xor (A(117) and B(9)) xor (A(118) and B(8)) xor (A(119) and B(7)) xor (A(120) and B(6)) xor (A(121) and B(5)) xor (A(122) and B(4)) xor (A(123) and B(3)) xor (A(124) and B(2)) xor (A(125) and B(1)) xor (A(126) and B(0)) xor (A(119) and B(127)) xor (A(120) and B(126)) xor (A(121) and B(125)) xor (A(122) and B(124)) xor (A(123) and B(123)) xor (A(124) and B(122)) xor (A(125) and B(121)) xor (A(126) and B(120)) xor (A(124) and B(127)) xor (A(125) and B(126)) xor (A(126) and B(125)) xor (A(125) and B(127)) xor (A(126) and B(126)) xor (A(126) and B(127));
    C(127) <= (A(0) and B(127)) xor (A(1) and B(126)) xor (A(2) and B(125)) xor (A(3) and B(124)) xor (A(4) and B(123)) xor (A(5) and B(122)) xor (A(6) and B(121)) xor (A(7) and B(120)) xor (A(8) and B(119)) xor (A(9) and B(118)) xor (A(10) and B(117)) xor (A(11) and B(116)) xor (A(12) and B(115)) xor (A(13) and B(114)) xor (A(14) and B(113)) xor (A(15) and B(112)) xor (A(16) and B(111)) xor (A(17) and B(110)) xor (A(18) and B(109)) xor (A(19) and B(108)) xor (A(20) and B(107)) xor (A(21) and B(106)) xor (A(23) and B(105)) xor (A(23) and B(104)) xor (A(24) and B(103)) xor (A(25) and B(102)) xor (A(26) and B(101)) xor (A(27) and B(100)) xor (A(28) and B(99)) xor (A(29) and B(98)) xor (A(30) and B(97)) xor (A(31) and B(96)) xor (A(32) and B(95)) xor (A(33) and B(94)) xor (A(34) and B(93)) xor (A(35) and B(92)) xor (A(36) and B(91)) xor (A(37) and B(90)) xor (A(38) and B(89)) xor (A(39) and B(88)) xor (A(40) and B(87)) xor (A(41) and B(86)) xor (A(42) and B(85)) xor (A(43) and B(84)) xor (A(44) and B(83)) xor (A(45) and B(82)) xor (A(46) and B(81)) xor (A(47) and B(80)) xor (A(48) and B(79)) xor (A(49) and B(78)) xor (A(50) and B(77)) xor (A(51) and B(76)) xor (A(52) and B(75)) xor (A(53) and B(74)) xor (A(54) and B(73)) xor (A(55) and B(72)) xor (A(56) and B(71)) xor (A(57) and B(70)) xor (A(58) and B(69)) xor (A(59) and B(68)) xor (A(60) and B(67)) xor (A(61) and B(66)) xor (A(62) and B(65)) xor (A(63) and B(64)) xor (A(64) and B(63)) xor (A(65) and B(62)) xor (A(66) and B(61)) xor (A(67) and B(60)) xor (A(68) and B(59)) xor (A(69) and B(58)) xor (A(70) and B(57)) xor (A(71) and B(56)) xor (A(72) and B(55)) xor (A(73) and B(54)) xor (A(74) and B(53)) xor (A(75) and B(52)) xor (A(76) and B(51)) xor (A(77) and B(50)) xor (A(78) and B(49)) xor (A(79) and B(48)) xor (A(80) and B(47)) xor (A(81) and B(46)) xor (A(82) and B(45)) xor (A(83) and B(44)) xor (A(84) and B(43)) xor (A(85) and B(42)) xor (A(86) and B(41)) xor (A(87) and B(40)) xor (A(88) and B(39)) xor (A(89) and B(38)) xor (A(90) and B(37)) xor (A(91) and B(36)) xor (A(92) and B(35)) xor (A(93) and B(34)) xor (A(94) and B(33)) xor (A(95) and B(32)) xor (A(96) and B(31)) xor (A(97) and B(30)) xor (A(98) and B(29)) xor (A(99) and B(28)) xor (A(100) and B(27)) xor (A(101) and B(26)) xor (A(102) and B(25)) xor (A(103) and B(24)) xor (A(104) and B(23)) xor (A(105) and B(23)) xor (A(106) and B(21)) xor (A(107) and B(20)) xor (A(108) and B(19)) xor (A(109) and B(18)) xor (A(110) and B(17)) xor (A(111) and B(16)) xor (A(112) and B(15)) xor (A(113) and B(14)) xor (A(114) and B(13)) xor (A(115) and B(12)) xor (A(116) and B(11)) xor (A(117) and B(10)) xor (A(118) and B(9)) xor (A(119) and B(8)) xor (A(120) and B(7)) xor (A(121) and B(6)) xor (A(122) and B(5)) xor (A(123) and B(4)) xor (A(124) and B(3)) xor (A(125) and B(2)) xor (A(126) and B(1)) xor (A(127) and B(0)) xor (A(120) and B(127)) xor (A(121) and B(126)) xor (A(122) and B(125)) xor (A(123) and B(124)) xor (A(124) and B(123)) xor (A(125) and B(122)) xor (A(126) and B(121)) xor (A(125) and B(127)) xor (A(126) and B(126)) xor (A(126) and B(127));

	PROCESS (clk)
	BEGIN
		IF rising_edge(clk) THEN
			IF (in_val = '1') THEN
				out_product <= C;
				out_val <= '1';
			ELSE
				out_val <= '0';
			END IF;
		END IF;
	END PROCESS;


END ARCHITECTURE;